module result_text_setter(clk, score, inresult, main_difficulty, x_pointer, y_pointer, result_text);
   input inresult;
	input [3:0] main_difficulty;
   input clk;
   input [7:0] x_pointer;
	input [6:0] y_pointer;
	input [12:0] score;
	output reg result_text; // check if the pixel is the menu's text.
	
	reg [3:0] units_digit_score;
	reg [3:0] tens_digit_score;
	reg [3:0] hundreds_digit_score;

	always@(posedge clk)begin
		units_digit_score <= score % 10;
	   tens_digit_score <= ((score - (score % 10)) / 10) % 10;
		hundreds_digit_score <= score / 100;
	end

	//menu's normal text
	always@(posedge clk)
	begin
		if (inresult)
			 begin
			 if (main_texts)
				 result_text <= 1'b1;
			 else
				 result_text <= 1'b0;
			 end
	end

	// wires for result texts
	wire main_texts = (x_pointer == 20 && y_pointer == 28)
||(x_pointer == 21 && y_pointer == 28)
||(x_pointer == 22 && y_pointer == 28)
||(x_pointer == 23 && y_pointer == 28)
||(x_pointer == 24 && y_pointer == 28)
||(x_pointer == 25 && y_pointer == 28)
||(x_pointer == 26 && y_pointer == 28)
||(x_pointer == 27 && y_pointer == 28)
||(x_pointer == 28 && y_pointer == 28)
||(x_pointer == 29 && y_pointer == 28)
||(x_pointer == 30 && y_pointer == 28)
||(x_pointer == 31 && y_pointer == 28)
||(x_pointer == 39 && y_pointer == 28)
||(x_pointer == 40 && y_pointer == 28)
||(x_pointer == 41 && y_pointer == 28)
||(x_pointer == 49 && y_pointer == 28)
||(x_pointer == 50 && y_pointer == 28)
||(x_pointer == 51 && y_pointer == 28)
||(x_pointer == 60 && y_pointer == 28)
||(x_pointer == 61 && y_pointer == 28)
||(x_pointer == 62 && y_pointer == 28)
||(x_pointer == 67 && y_pointer == 28)
||(x_pointer == 68 && y_pointer == 28)
||(x_pointer == 69 && y_pointer == 28)
||(x_pointer == 70 && y_pointer == 28)
||(x_pointer == 71 && y_pointer == 28)
||(x_pointer == 72 && y_pointer == 28)
||(x_pointer == 73 && y_pointer == 28)
||(x_pointer == 74 && y_pointer == 28)
||(x_pointer == 75 && y_pointer == 28)
||(x_pointer == 76 && y_pointer == 28)
||(x_pointer == 87 && y_pointer == 28)
||(x_pointer == 88 && y_pointer == 28)
||(x_pointer == 89 && y_pointer == 28)
||(x_pointer == 90 && y_pointer == 28)
||(x_pointer == 91 && y_pointer == 28)
||(x_pointer == 92 && y_pointer == 28)
||(x_pointer == 93 && y_pointer == 28)
||(x_pointer == 94 && y_pointer == 28)
||(x_pointer == 95 && y_pointer == 28)
||(x_pointer == 96 && y_pointer == 28)
||(x_pointer == 97 && y_pointer == 28)
||(x_pointer == 98 && y_pointer == 28)
||(x_pointer == 102 && y_pointer == 28)
||(x_pointer == 103 && y_pointer == 28)
||(x_pointer == 104 && y_pointer == 28)
||(x_pointer == 111 && y_pointer == 28)
||(x_pointer == 112 && y_pointer == 28)
||(x_pointer == 113 && y_pointer == 28)
||(x_pointer == 117 && y_pointer == 28)
||(x_pointer == 118 && y_pointer == 28)
||(x_pointer == 119 && y_pointer == 28)
||(x_pointer == 120 && y_pointer == 28)
||(x_pointer == 121 && y_pointer == 28)
||(x_pointer == 122 && y_pointer == 28)
||(x_pointer == 123 && y_pointer == 28)
||(x_pointer == 124 && y_pointer == 28)
||(x_pointer == 125 && y_pointer == 28)
||(x_pointer == 126 && y_pointer == 28)
||(x_pointer == 130 && y_pointer == 28)
||(x_pointer == 131 && y_pointer == 28)
||(x_pointer == 132 && y_pointer == 28)
||(x_pointer == 133 && y_pointer == 28)
||(x_pointer == 134 && y_pointer == 28)
||(x_pointer == 135 && y_pointer == 28)
||(x_pointer == 136 && y_pointer == 28)
||(x_pointer == 137 && y_pointer == 28)
||(x_pointer == 138 && y_pointer == 28)
||(x_pointer == 139 && y_pointer == 28)
||(x_pointer == 140 && y_pointer == 28)
||(x_pointer == 141 && y_pointer == 28)
||(x_pointer == 20 && y_pointer == 29)
||(x_pointer == 21 && y_pointer == 29)
||(x_pointer == 22 && y_pointer == 29)
||(x_pointer == 23 && y_pointer == 29)
||(x_pointer == 24 && y_pointer == 29)
||(x_pointer == 25 && y_pointer == 29)
||(x_pointer == 26 && y_pointer == 29)
||(x_pointer == 27 && y_pointer == 29)
||(x_pointer == 28 && y_pointer == 29)
||(x_pointer == 29 && y_pointer == 29)
||(x_pointer == 30 && y_pointer == 29)
||(x_pointer == 31 && y_pointer == 29)
||(x_pointer == 39 && y_pointer == 29)
||(x_pointer == 40 && y_pointer == 29)
||(x_pointer == 41 && y_pointer == 29)
||(x_pointer == 49 && y_pointer == 29)
||(x_pointer == 50 && y_pointer == 29)
||(x_pointer == 51 && y_pointer == 29)
||(x_pointer == 60 && y_pointer == 29)
||(x_pointer == 61 && y_pointer == 29)
||(x_pointer == 62 && y_pointer == 29)
||(x_pointer == 67 && y_pointer == 29)
||(x_pointer == 68 && y_pointer == 29)
||(x_pointer == 69 && y_pointer == 29)
||(x_pointer == 70 && y_pointer == 29)
||(x_pointer == 71 && y_pointer == 29)
||(x_pointer == 72 && y_pointer == 29)
||(x_pointer == 73 && y_pointer == 29)
||(x_pointer == 74 && y_pointer == 29)
||(x_pointer == 75 && y_pointer == 29)
||(x_pointer == 76 && y_pointer == 29)
||(x_pointer == 87 && y_pointer == 29)
||(x_pointer == 88 && y_pointer == 29)
||(x_pointer == 89 && y_pointer == 29)
||(x_pointer == 90 && y_pointer == 29)
||(x_pointer == 91 && y_pointer == 29)
||(x_pointer == 92 && y_pointer == 29)
||(x_pointer == 93 && y_pointer == 29)
||(x_pointer == 94 && y_pointer == 29)
||(x_pointer == 95 && y_pointer == 29)
||(x_pointer == 96 && y_pointer == 29)
||(x_pointer == 97 && y_pointer == 29)
||(x_pointer == 98 && y_pointer == 29)
||(x_pointer == 102 && y_pointer == 29)
||(x_pointer == 103 && y_pointer == 29)
||(x_pointer == 104 && y_pointer == 29)
||(x_pointer == 111 && y_pointer == 29)
||(x_pointer == 112 && y_pointer == 29)
||(x_pointer == 113 && y_pointer == 29)
||(x_pointer == 117 && y_pointer == 29)
||(x_pointer == 118 && y_pointer == 29)
||(x_pointer == 119 && y_pointer == 29)
||(x_pointer == 120 && y_pointer == 29)
||(x_pointer == 121 && y_pointer == 29)
||(x_pointer == 122 && y_pointer == 29)
||(x_pointer == 123 && y_pointer == 29)
||(x_pointer == 124 && y_pointer == 29)
||(x_pointer == 125 && y_pointer == 29)
||(x_pointer == 126 && y_pointer == 29)
||(x_pointer == 130 && y_pointer == 29)
||(x_pointer == 131 && y_pointer == 29)
||(x_pointer == 132 && y_pointer == 29)
||(x_pointer == 133 && y_pointer == 29)
||(x_pointer == 134 && y_pointer == 29)
||(x_pointer == 135 && y_pointer == 29)
||(x_pointer == 136 && y_pointer == 29)
||(x_pointer == 137 && y_pointer == 29)
||(x_pointer == 138 && y_pointer == 29)
||(x_pointer == 139 && y_pointer == 29)
||(x_pointer == 140 && y_pointer == 29)
||(x_pointer == 141 && y_pointer == 29)
||(x_pointer == 20 && y_pointer == 30)
||(x_pointer == 21 && y_pointer == 30)
||(x_pointer == 22 && y_pointer == 30)
||(x_pointer == 28 && y_pointer == 30)
||(x_pointer == 29 && y_pointer == 30)
||(x_pointer == 30 && y_pointer == 30)
||(x_pointer == 31 && y_pointer == 30)
||(x_pointer == 38 && y_pointer == 30)
||(x_pointer == 39 && y_pointer == 30)
||(x_pointer == 40 && y_pointer == 30)
||(x_pointer == 41 && y_pointer == 30)
||(x_pointer == 42 && y_pointer == 30)
||(x_pointer == 49 && y_pointer == 30)
||(x_pointer == 50 && y_pointer == 30)
||(x_pointer == 51 && y_pointer == 30)
||(x_pointer == 52 && y_pointer == 30)
||(x_pointer == 59 && y_pointer == 30)
||(x_pointer == 60 && y_pointer == 30)
||(x_pointer == 61 && y_pointer == 30)
||(x_pointer == 62 && y_pointer == 30)
||(x_pointer == 67 && y_pointer == 30)
||(x_pointer == 68 && y_pointer == 30)
||(x_pointer == 69 && y_pointer == 30)
||(x_pointer == 87 && y_pointer == 30)
||(x_pointer == 88 && y_pointer == 30)
||(x_pointer == 89 && y_pointer == 30)
||(x_pointer == 96 && y_pointer == 30)
||(x_pointer == 97 && y_pointer == 30)
||(x_pointer == 98 && y_pointer == 30)
||(x_pointer == 102 && y_pointer == 30)
||(x_pointer == 103 && y_pointer == 30)
||(x_pointer == 104 && y_pointer == 30)
||(x_pointer == 111 && y_pointer == 30)
||(x_pointer == 112 && y_pointer == 30)
||(x_pointer == 113 && y_pointer == 30)
||(x_pointer == 117 && y_pointer == 30)
||(x_pointer == 118 && y_pointer == 30)
||(x_pointer == 119 && y_pointer == 30)
||(x_pointer == 130 && y_pointer == 30)
||(x_pointer == 131 && y_pointer == 30)
||(x_pointer == 132 && y_pointer == 30)
||(x_pointer == 138 && y_pointer == 30)
||(x_pointer == 139 && y_pointer == 30)
||(x_pointer == 140 && y_pointer == 30)
||(x_pointer == 141 && y_pointer == 30)
||(x_pointer == 20 && y_pointer == 31)
||(x_pointer == 21 && y_pointer == 31)
||(x_pointer == 22 && y_pointer == 31)
||(x_pointer == 28 && y_pointer == 31)
||(x_pointer == 29 && y_pointer == 31)
||(x_pointer == 30 && y_pointer == 31)
||(x_pointer == 31 && y_pointer == 31)
||(x_pointer == 38 && y_pointer == 31)
||(x_pointer == 39 && y_pointer == 31)
||(x_pointer == 40 && y_pointer == 31)
||(x_pointer == 41 && y_pointer == 31)
||(x_pointer == 42 && y_pointer == 31)
||(x_pointer == 49 && y_pointer == 31)
||(x_pointer == 50 && y_pointer == 31)
||(x_pointer == 51 && y_pointer == 31)
||(x_pointer == 52 && y_pointer == 31)
||(x_pointer == 59 && y_pointer == 31)
||(x_pointer == 60 && y_pointer == 31)
||(x_pointer == 61 && y_pointer == 31)
||(x_pointer == 62 && y_pointer == 31)
||(x_pointer == 67 && y_pointer == 31)
||(x_pointer == 68 && y_pointer == 31)
||(x_pointer == 69 && y_pointer == 31)
||(x_pointer == 87 && y_pointer == 31)
||(x_pointer == 88 && y_pointer == 31)
||(x_pointer == 89 && y_pointer == 31)
||(x_pointer == 96 && y_pointer == 31)
||(x_pointer == 97 && y_pointer == 31)
||(x_pointer == 98 && y_pointer == 31)
||(x_pointer == 102 && y_pointer == 31)
||(x_pointer == 103 && y_pointer == 31)
||(x_pointer == 104 && y_pointer == 31)
||(x_pointer == 105 && y_pointer == 31)
||(x_pointer == 110 && y_pointer == 31)
||(x_pointer == 111 && y_pointer == 31)
||(x_pointer == 112 && y_pointer == 31)
||(x_pointer == 113 && y_pointer == 31)
||(x_pointer == 117 && y_pointer == 31)
||(x_pointer == 118 && y_pointer == 31)
||(x_pointer == 119 && y_pointer == 31)
||(x_pointer == 130 && y_pointer == 31)
||(x_pointer == 131 && y_pointer == 31)
||(x_pointer == 132 && y_pointer == 31)
||(x_pointer == 138 && y_pointer == 31)
||(x_pointer == 139 && y_pointer == 31)
||(x_pointer == 140 && y_pointer == 31)
||(x_pointer == 141 && y_pointer == 31)
||(x_pointer == 20 && y_pointer == 32)
||(x_pointer == 21 && y_pointer == 32)
||(x_pointer == 22 && y_pointer == 32)
||(x_pointer == 28 && y_pointer == 32)
||(x_pointer == 29 && y_pointer == 32)
||(x_pointer == 30 && y_pointer == 32)
||(x_pointer == 31 && y_pointer == 32)
||(x_pointer == 38 && y_pointer == 32)
||(x_pointer == 39 && y_pointer == 32)
||(x_pointer == 40 && y_pointer == 32)
||(x_pointer == 41 && y_pointer == 32)
||(x_pointer == 42 && y_pointer == 32)
||(x_pointer == 49 && y_pointer == 32)
||(x_pointer == 50 && y_pointer == 32)
||(x_pointer == 51 && y_pointer == 32)
||(x_pointer == 52 && y_pointer == 32)
||(x_pointer == 59 && y_pointer == 32)
||(x_pointer == 60 && y_pointer == 32)
||(x_pointer == 61 && y_pointer == 32)
||(x_pointer == 62 && y_pointer == 32)
||(x_pointer == 67 && y_pointer == 32)
||(x_pointer == 68 && y_pointer == 32)
||(x_pointer == 69 && y_pointer == 32)
||(x_pointer == 87 && y_pointer == 32)
||(x_pointer == 88 && y_pointer == 32)
||(x_pointer == 89 && y_pointer == 32)
||(x_pointer == 96 && y_pointer == 32)
||(x_pointer == 97 && y_pointer == 32)
||(x_pointer == 98 && y_pointer == 32)
||(x_pointer == 103 && y_pointer == 32)
||(x_pointer == 104 && y_pointer == 32)
||(x_pointer == 105 && y_pointer == 32)
||(x_pointer == 110 && y_pointer == 32)
||(x_pointer == 111 && y_pointer == 32)
||(x_pointer == 112 && y_pointer == 32)
||(x_pointer == 117 && y_pointer == 32)
||(x_pointer == 118 && y_pointer == 32)
||(x_pointer == 119 && y_pointer == 32)
||(x_pointer == 130 && y_pointer == 32)
||(x_pointer == 131 && y_pointer == 32)
||(x_pointer == 132 && y_pointer == 32)
||(x_pointer == 138 && y_pointer == 32)
||(x_pointer == 139 && y_pointer == 32)
||(x_pointer == 140 && y_pointer == 32)
||(x_pointer == 141 && y_pointer == 32)
||(x_pointer == 20 && y_pointer == 33)
||(x_pointer == 21 && y_pointer == 33)
||(x_pointer == 22 && y_pointer == 33)
||(x_pointer == 28 && y_pointer == 33)
||(x_pointer == 29 && y_pointer == 33)
||(x_pointer == 30 && y_pointer == 33)
||(x_pointer == 31 && y_pointer == 33)
||(x_pointer == 38 && y_pointer == 33)
||(x_pointer == 39 && y_pointer == 33)
||(x_pointer == 40 && y_pointer == 33)
||(x_pointer == 41 && y_pointer == 33)
||(x_pointer == 42 && y_pointer == 33)
||(x_pointer == 49 && y_pointer == 33)
||(x_pointer == 50 && y_pointer == 33)
||(x_pointer == 51 && y_pointer == 33)
||(x_pointer == 52 && y_pointer == 33)
||(x_pointer == 53 && y_pointer == 33)
||(x_pointer == 58 && y_pointer == 33)
||(x_pointer == 59 && y_pointer == 33)
||(x_pointer == 60 && y_pointer == 33)
||(x_pointer == 61 && y_pointer == 33)
||(x_pointer == 62 && y_pointer == 33)
||(x_pointer == 67 && y_pointer == 33)
||(x_pointer == 68 && y_pointer == 33)
||(x_pointer == 69 && y_pointer == 33)
||(x_pointer == 87 && y_pointer == 33)
||(x_pointer == 88 && y_pointer == 33)
||(x_pointer == 89 && y_pointer == 33)
||(x_pointer == 96 && y_pointer == 33)
||(x_pointer == 97 && y_pointer == 33)
||(x_pointer == 98 && y_pointer == 33)
||(x_pointer == 103 && y_pointer == 33)
||(x_pointer == 104 && y_pointer == 33)
||(x_pointer == 105 && y_pointer == 33)
||(x_pointer == 110 && y_pointer == 33)
||(x_pointer == 111 && y_pointer == 33)
||(x_pointer == 112 && y_pointer == 33)
||(x_pointer == 117 && y_pointer == 33)
||(x_pointer == 118 && y_pointer == 33)
||(x_pointer == 119 && y_pointer == 33)
||(x_pointer == 130 && y_pointer == 33)
||(x_pointer == 131 && y_pointer == 33)
||(x_pointer == 132 && y_pointer == 33)
||(x_pointer == 138 && y_pointer == 33)
||(x_pointer == 139 && y_pointer == 33)
||(x_pointer == 140 && y_pointer == 33)
||(x_pointer == 141 && y_pointer == 33)
||(x_pointer == 20 && y_pointer == 34)
||(x_pointer == 21 && y_pointer == 34)
||(x_pointer == 22 && y_pointer == 34)
||(x_pointer == 28 && y_pointer == 34)
||(x_pointer == 29 && y_pointer == 34)
||(x_pointer == 30 && y_pointer == 34)
||(x_pointer == 31 && y_pointer == 34)
||(x_pointer == 37 && y_pointer == 34)
||(x_pointer == 38 && y_pointer == 34)
||(x_pointer == 39 && y_pointer == 34)
||(x_pointer == 40 && y_pointer == 34)
||(x_pointer == 41 && y_pointer == 34)
||(x_pointer == 42 && y_pointer == 34)
||(x_pointer == 43 && y_pointer == 34)
||(x_pointer == 49 && y_pointer == 34)
||(x_pointer == 50 && y_pointer == 34)
||(x_pointer == 51 && y_pointer == 34)
||(x_pointer == 52 && y_pointer == 34)
||(x_pointer == 53 && y_pointer == 34)
||(x_pointer == 58 && y_pointer == 34)
||(x_pointer == 59 && y_pointer == 34)
||(x_pointer == 60 && y_pointer == 34)
||(x_pointer == 61 && y_pointer == 34)
||(x_pointer == 62 && y_pointer == 34)
||(x_pointer == 67 && y_pointer == 34)
||(x_pointer == 68 && y_pointer == 34)
||(x_pointer == 69 && y_pointer == 34)
||(x_pointer == 87 && y_pointer == 34)
||(x_pointer == 88 && y_pointer == 34)
||(x_pointer == 89 && y_pointer == 34)
||(x_pointer == 96 && y_pointer == 34)
||(x_pointer == 97 && y_pointer == 34)
||(x_pointer == 98 && y_pointer == 34)
||(x_pointer == 103 && y_pointer == 34)
||(x_pointer == 104 && y_pointer == 34)
||(x_pointer == 105 && y_pointer == 34)
||(x_pointer == 110 && y_pointer == 34)
||(x_pointer == 111 && y_pointer == 34)
||(x_pointer == 112 && y_pointer == 34)
||(x_pointer == 117 && y_pointer == 34)
||(x_pointer == 118 && y_pointer == 34)
||(x_pointer == 119 && y_pointer == 34)
||(x_pointer == 130 && y_pointer == 34)
||(x_pointer == 131 && y_pointer == 34)
||(x_pointer == 132 && y_pointer == 34)
||(x_pointer == 138 && y_pointer == 34)
||(x_pointer == 139 && y_pointer == 34)
||(x_pointer == 140 && y_pointer == 34)
||(x_pointer == 141 && y_pointer == 34)
||(x_pointer == 20 && y_pointer == 35)
||(x_pointer == 21 && y_pointer == 35)
||(x_pointer == 22 && y_pointer == 35)
||(x_pointer == 37 && y_pointer == 35)
||(x_pointer == 38 && y_pointer == 35)
||(x_pointer == 39 && y_pointer == 35)
||(x_pointer == 40 && y_pointer == 35)
||(x_pointer == 41 && y_pointer == 35)
||(x_pointer == 42 && y_pointer == 35)
||(x_pointer == 43 && y_pointer == 35)
||(x_pointer == 49 && y_pointer == 35)
||(x_pointer == 50 && y_pointer == 35)
||(x_pointer == 51 && y_pointer == 35)
||(x_pointer == 52 && y_pointer == 35)
||(x_pointer == 53 && y_pointer == 35)
||(x_pointer == 58 && y_pointer == 35)
||(x_pointer == 59 && y_pointer == 35)
||(x_pointer == 60 && y_pointer == 35)
||(x_pointer == 61 && y_pointer == 35)
||(x_pointer == 62 && y_pointer == 35)
||(x_pointer == 67 && y_pointer == 35)
||(x_pointer == 68 && y_pointer == 35)
||(x_pointer == 69 && y_pointer == 35)
||(x_pointer == 87 && y_pointer == 35)
||(x_pointer == 88 && y_pointer == 35)
||(x_pointer == 89 && y_pointer == 35)
||(x_pointer == 96 && y_pointer == 35)
||(x_pointer == 97 && y_pointer == 35)
||(x_pointer == 98 && y_pointer == 35)
||(x_pointer == 103 && y_pointer == 35)
||(x_pointer == 104 && y_pointer == 35)
||(x_pointer == 105 && y_pointer == 35)
||(x_pointer == 110 && y_pointer == 35)
||(x_pointer == 111 && y_pointer == 35)
||(x_pointer == 112 && y_pointer == 35)
||(x_pointer == 117 && y_pointer == 35)
||(x_pointer == 118 && y_pointer == 35)
||(x_pointer == 119 && y_pointer == 35)
||(x_pointer == 130 && y_pointer == 35)
||(x_pointer == 131 && y_pointer == 35)
||(x_pointer == 132 && y_pointer == 35)
||(x_pointer == 138 && y_pointer == 35)
||(x_pointer == 139 && y_pointer == 35)
||(x_pointer == 140 && y_pointer == 35)
||(x_pointer == 141 && y_pointer == 35)
||(x_pointer == 20 && y_pointer == 36)
||(x_pointer == 21 && y_pointer == 36)
||(x_pointer == 22 && y_pointer == 36)
||(x_pointer == 37 && y_pointer == 36)
||(x_pointer == 38 && y_pointer == 36)
||(x_pointer == 39 && y_pointer == 36)
||(x_pointer == 41 && y_pointer == 36)
||(x_pointer == 42 && y_pointer == 36)
||(x_pointer == 43 && y_pointer == 36)
||(x_pointer == 49 && y_pointer == 36)
||(x_pointer == 50 && y_pointer == 36)
||(x_pointer == 51 && y_pointer == 36)
||(x_pointer == 52 && y_pointer == 36)
||(x_pointer == 53 && y_pointer == 36)
||(x_pointer == 54 && y_pointer == 36)
||(x_pointer == 57 && y_pointer == 36)
||(x_pointer == 58 && y_pointer == 36)
||(x_pointer == 59 && y_pointer == 36)
||(x_pointer == 60 && y_pointer == 36)
||(x_pointer == 61 && y_pointer == 36)
||(x_pointer == 62 && y_pointer == 36)
||(x_pointer == 67 && y_pointer == 36)
||(x_pointer == 68 && y_pointer == 36)
||(x_pointer == 69 && y_pointer == 36)
||(x_pointer == 87 && y_pointer == 36)
||(x_pointer == 88 && y_pointer == 36)
||(x_pointer == 89 && y_pointer == 36)
||(x_pointer == 96 && y_pointer == 36)
||(x_pointer == 97 && y_pointer == 36)
||(x_pointer == 98 && y_pointer == 36)
||(x_pointer == 104 && y_pointer == 36)
||(x_pointer == 105 && y_pointer == 36)
||(x_pointer == 106 && y_pointer == 36)
||(x_pointer == 109 && y_pointer == 36)
||(x_pointer == 110 && y_pointer == 36)
||(x_pointer == 111 && y_pointer == 36)
||(x_pointer == 112 && y_pointer == 36)
||(x_pointer == 117 && y_pointer == 36)
||(x_pointer == 118 && y_pointer == 36)
||(x_pointer == 119 && y_pointer == 36)
||(x_pointer == 130 && y_pointer == 36)
||(x_pointer == 131 && y_pointer == 36)
||(x_pointer == 132 && y_pointer == 36)
||(x_pointer == 138 && y_pointer == 36)
||(x_pointer == 139 && y_pointer == 36)
||(x_pointer == 140 && y_pointer == 36)
||(x_pointer == 141 && y_pointer == 36)
||(x_pointer == 20 && y_pointer == 37)
||(x_pointer == 21 && y_pointer == 37)
||(x_pointer == 22 && y_pointer == 37)
||(x_pointer == 37 && y_pointer == 37)
||(x_pointer == 38 && y_pointer == 37)
||(x_pointer == 39 && y_pointer == 37)
||(x_pointer == 41 && y_pointer == 37)
||(x_pointer == 42 && y_pointer == 37)
||(x_pointer == 43 && y_pointer == 37)
||(x_pointer == 49 && y_pointer == 37)
||(x_pointer == 50 && y_pointer == 37)
||(x_pointer == 51 && y_pointer == 37)
||(x_pointer == 52 && y_pointer == 37)
||(x_pointer == 53 && y_pointer == 37)
||(x_pointer == 54 && y_pointer == 37)
||(x_pointer == 57 && y_pointer == 37)
||(x_pointer == 58 && y_pointer == 37)
||(x_pointer == 59 && y_pointer == 37)
||(x_pointer == 60 && y_pointer == 37)
||(x_pointer == 61 && y_pointer == 37)
||(x_pointer == 62 && y_pointer == 37)
||(x_pointer == 67 && y_pointer == 37)
||(x_pointer == 68 && y_pointer == 37)
||(x_pointer == 69 && y_pointer == 37)
||(x_pointer == 70 && y_pointer == 37)
||(x_pointer == 71 && y_pointer == 37)
||(x_pointer == 72 && y_pointer == 37)
||(x_pointer == 73 && y_pointer == 37)
||(x_pointer == 74 && y_pointer == 37)
||(x_pointer == 75 && y_pointer == 37)
||(x_pointer == 87 && y_pointer == 37)
||(x_pointer == 88 && y_pointer == 37)
||(x_pointer == 89 && y_pointer == 37)
||(x_pointer == 96 && y_pointer == 37)
||(x_pointer == 97 && y_pointer == 37)
||(x_pointer == 98 && y_pointer == 37)
||(x_pointer == 104 && y_pointer == 37)
||(x_pointer == 105 && y_pointer == 37)
||(x_pointer == 106 && y_pointer == 37)
||(x_pointer == 109 && y_pointer == 37)
||(x_pointer == 110 && y_pointer == 37)
||(x_pointer == 111 && y_pointer == 37)
||(x_pointer == 117 && y_pointer == 37)
||(x_pointer == 118 && y_pointer == 37)
||(x_pointer == 119 && y_pointer == 37)
||(x_pointer == 120 && y_pointer == 37)
||(x_pointer == 121 && y_pointer == 37)
||(x_pointer == 122 && y_pointer == 37)
||(x_pointer == 123 && y_pointer == 37)
||(x_pointer == 124 && y_pointer == 37)
||(x_pointer == 125 && y_pointer == 37)
||(x_pointer == 130 && y_pointer == 37)
||(x_pointer == 131 && y_pointer == 37)
||(x_pointer == 132 && y_pointer == 37)
||(x_pointer == 134 && y_pointer == 37)
||(x_pointer == 135 && y_pointer == 37)
||(x_pointer == 136 && y_pointer == 37)
||(x_pointer == 137 && y_pointer == 37)
||(x_pointer == 138 && y_pointer == 37)
||(x_pointer == 139 && y_pointer == 37)
||(x_pointer == 140 && y_pointer == 37)
||(x_pointer == 141 && y_pointer == 37)
||(x_pointer == 20 && y_pointer == 38)
||(x_pointer == 21 && y_pointer == 38)
||(x_pointer == 22 && y_pointer == 38)
||(x_pointer == 25 && y_pointer == 38)
||(x_pointer == 26 && y_pointer == 38)
||(x_pointer == 27 && y_pointer == 38)
||(x_pointer == 28 && y_pointer == 38)
||(x_pointer == 29 && y_pointer == 38)
||(x_pointer == 30 && y_pointer == 38)
||(x_pointer == 31 && y_pointer == 38)
||(x_pointer == 36 && y_pointer == 38)
||(x_pointer == 37 && y_pointer == 38)
||(x_pointer == 38 && y_pointer == 38)
||(x_pointer == 39 && y_pointer == 38)
||(x_pointer == 41 && y_pointer == 38)
||(x_pointer == 42 && y_pointer == 38)
||(x_pointer == 43 && y_pointer == 38)
||(x_pointer == 44 && y_pointer == 38)
||(x_pointer == 49 && y_pointer == 38)
||(x_pointer == 50 && y_pointer == 38)
||(x_pointer == 51 && y_pointer == 38)
||(x_pointer == 52 && y_pointer == 38)
||(x_pointer == 53 && y_pointer == 38)
||(x_pointer == 54 && y_pointer == 38)
||(x_pointer == 57 && y_pointer == 38)
||(x_pointer == 58 && y_pointer == 38)
||(x_pointer == 59 && y_pointer == 38)
||(x_pointer == 60 && y_pointer == 38)
||(x_pointer == 61 && y_pointer == 38)
||(x_pointer == 62 && y_pointer == 38)
||(x_pointer == 67 && y_pointer == 38)
||(x_pointer == 68 && y_pointer == 38)
||(x_pointer == 69 && y_pointer == 38)
||(x_pointer == 70 && y_pointer == 38)
||(x_pointer == 71 && y_pointer == 38)
||(x_pointer == 72 && y_pointer == 38)
||(x_pointer == 73 && y_pointer == 38)
||(x_pointer == 74 && y_pointer == 38)
||(x_pointer == 75 && y_pointer == 38)
||(x_pointer == 87 && y_pointer == 38)
||(x_pointer == 88 && y_pointer == 38)
||(x_pointer == 89 && y_pointer == 38)
||(x_pointer == 96 && y_pointer == 38)
||(x_pointer == 97 && y_pointer == 38)
||(x_pointer == 98 && y_pointer == 38)
||(x_pointer == 104 && y_pointer == 38)
||(x_pointer == 105 && y_pointer == 38)
||(x_pointer == 106 && y_pointer == 38)
||(x_pointer == 109 && y_pointer == 38)
||(x_pointer == 110 && y_pointer == 38)
||(x_pointer == 111 && y_pointer == 38)
||(x_pointer == 117 && y_pointer == 38)
||(x_pointer == 118 && y_pointer == 38)
||(x_pointer == 119 && y_pointer == 38)
||(x_pointer == 120 && y_pointer == 38)
||(x_pointer == 121 && y_pointer == 38)
||(x_pointer == 122 && y_pointer == 38)
||(x_pointer == 123 && y_pointer == 38)
||(x_pointer == 124 && y_pointer == 38)
||(x_pointer == 125 && y_pointer == 38)
||(x_pointer == 130 && y_pointer == 38)
||(x_pointer == 131 && y_pointer == 38)
||(x_pointer == 132 && y_pointer == 38)
||(x_pointer == 134 && y_pointer == 38)
||(x_pointer == 135 && y_pointer == 38)
||(x_pointer == 136 && y_pointer == 38)
||(x_pointer == 137 && y_pointer == 38)
||(x_pointer == 138 && y_pointer == 38)
||(x_pointer == 139 && y_pointer == 38)
||(x_pointer == 140 && y_pointer == 38)
||(x_pointer == 141 && y_pointer == 38)
||(x_pointer == 20 && y_pointer == 39)
||(x_pointer == 21 && y_pointer == 39)
||(x_pointer == 22 && y_pointer == 39)
||(x_pointer == 25 && y_pointer == 39)
||(x_pointer == 26 && y_pointer == 39)
||(x_pointer == 27 && y_pointer == 39)
||(x_pointer == 28 && y_pointer == 39)
||(x_pointer == 29 && y_pointer == 39)
||(x_pointer == 30 && y_pointer == 39)
||(x_pointer == 31 && y_pointer == 39)
||(x_pointer == 36 && y_pointer == 39)
||(x_pointer == 37 && y_pointer == 39)
||(x_pointer == 38 && y_pointer == 39)
||(x_pointer == 39 && y_pointer == 39)
||(x_pointer == 41 && y_pointer == 39)
||(x_pointer == 42 && y_pointer == 39)
||(x_pointer == 43 && y_pointer == 39)
||(x_pointer == 44 && y_pointer == 39)
||(x_pointer == 49 && y_pointer == 39)
||(x_pointer == 50 && y_pointer == 39)
||(x_pointer == 51 && y_pointer == 39)
||(x_pointer == 53 && y_pointer == 39)
||(x_pointer == 54 && y_pointer == 39)
||(x_pointer == 55 && y_pointer == 39)
||(x_pointer == 56 && y_pointer == 39)
||(x_pointer == 57 && y_pointer == 39)
||(x_pointer == 58 && y_pointer == 39)
||(x_pointer == 60 && y_pointer == 39)
||(x_pointer == 61 && y_pointer == 39)
||(x_pointer == 62 && y_pointer == 39)
||(x_pointer == 67 && y_pointer == 39)
||(x_pointer == 68 && y_pointer == 39)
||(x_pointer == 69 && y_pointer == 39)
||(x_pointer == 87 && y_pointer == 39)
||(x_pointer == 88 && y_pointer == 39)
||(x_pointer == 89 && y_pointer == 39)
||(x_pointer == 96 && y_pointer == 39)
||(x_pointer == 97 && y_pointer == 39)
||(x_pointer == 98 && y_pointer == 39)
||(x_pointer == 104 && y_pointer == 39)
||(x_pointer == 105 && y_pointer == 39)
||(x_pointer == 106 && y_pointer == 39)
||(x_pointer == 109 && y_pointer == 39)
||(x_pointer == 110 && y_pointer == 39)
||(x_pointer == 111 && y_pointer == 39)
||(x_pointer == 117 && y_pointer == 39)
||(x_pointer == 118 && y_pointer == 39)
||(x_pointer == 119 && y_pointer == 39)
||(x_pointer == 130 && y_pointer == 39)
||(x_pointer == 131 && y_pointer == 39)
||(x_pointer == 132 && y_pointer == 39)
||(x_pointer == 135 && y_pointer == 39)
||(x_pointer == 136 && y_pointer == 39)
||(x_pointer == 137 && y_pointer == 39)
||(x_pointer == 20 && y_pointer == 40)
||(x_pointer == 21 && y_pointer == 40)
||(x_pointer == 22 && y_pointer == 40)
||(x_pointer == 28 && y_pointer == 40)
||(x_pointer == 29 && y_pointer == 40)
||(x_pointer == 30 && y_pointer == 40)
||(x_pointer == 31 && y_pointer == 40)
||(x_pointer == 36 && y_pointer == 40)
||(x_pointer == 37 && y_pointer == 40)
||(x_pointer == 38 && y_pointer == 40)
||(x_pointer == 42 && y_pointer == 40)
||(x_pointer == 43 && y_pointer == 40)
||(x_pointer == 44 && y_pointer == 40)
||(x_pointer == 49 && y_pointer == 40)
||(x_pointer == 50 && y_pointer == 40)
||(x_pointer == 51 && y_pointer == 40)
||(x_pointer == 53 && y_pointer == 40)
||(x_pointer == 54 && y_pointer == 40)
||(x_pointer == 55 && y_pointer == 40)
||(x_pointer == 56 && y_pointer == 40)
||(x_pointer == 57 && y_pointer == 40)
||(x_pointer == 58 && y_pointer == 40)
||(x_pointer == 60 && y_pointer == 40)
||(x_pointer == 61 && y_pointer == 40)
||(x_pointer == 62 && y_pointer == 40)
||(x_pointer == 67 && y_pointer == 40)
||(x_pointer == 68 && y_pointer == 40)
||(x_pointer == 69 && y_pointer == 40)
||(x_pointer == 87 && y_pointer == 40)
||(x_pointer == 88 && y_pointer == 40)
||(x_pointer == 89 && y_pointer == 40)
||(x_pointer == 96 && y_pointer == 40)
||(x_pointer == 97 && y_pointer == 40)
||(x_pointer == 98 && y_pointer == 40)
||(x_pointer == 104 && y_pointer == 40)
||(x_pointer == 105 && y_pointer == 40)
||(x_pointer == 106 && y_pointer == 40)
||(x_pointer == 109 && y_pointer == 40)
||(x_pointer == 110 && y_pointer == 40)
||(x_pointer == 111 && y_pointer == 40)
||(x_pointer == 117 && y_pointer == 40)
||(x_pointer == 118 && y_pointer == 40)
||(x_pointer == 119 && y_pointer == 40)
||(x_pointer == 130 && y_pointer == 40)
||(x_pointer == 131 && y_pointer == 40)
||(x_pointer == 132 && y_pointer == 40)
||(x_pointer == 135 && y_pointer == 40)
||(x_pointer == 136 && y_pointer == 40)
||(x_pointer == 137 && y_pointer == 40)
||(x_pointer == 20 && y_pointer == 41)
||(x_pointer == 21 && y_pointer == 41)
||(x_pointer == 22 && y_pointer == 41)
||(x_pointer == 28 && y_pointer == 41)
||(x_pointer == 29 && y_pointer == 41)
||(x_pointer == 30 && y_pointer == 41)
||(x_pointer == 31 && y_pointer == 41)
||(x_pointer == 36 && y_pointer == 41)
||(x_pointer == 37 && y_pointer == 41)
||(x_pointer == 38 && y_pointer == 41)
||(x_pointer == 42 && y_pointer == 41)
||(x_pointer == 43 && y_pointer == 41)
||(x_pointer == 44 && y_pointer == 41)
||(x_pointer == 49 && y_pointer == 41)
||(x_pointer == 50 && y_pointer == 41)
||(x_pointer == 51 && y_pointer == 41)
||(x_pointer == 53 && y_pointer == 41)
||(x_pointer == 54 && y_pointer == 41)
||(x_pointer == 55 && y_pointer == 41)
||(x_pointer == 56 && y_pointer == 41)
||(x_pointer == 57 && y_pointer == 41)
||(x_pointer == 58 && y_pointer == 41)
||(x_pointer == 60 && y_pointer == 41)
||(x_pointer == 61 && y_pointer == 41)
||(x_pointer == 62 && y_pointer == 41)
||(x_pointer == 67 && y_pointer == 41)
||(x_pointer == 68 && y_pointer == 41)
||(x_pointer == 69 && y_pointer == 41)
||(x_pointer == 87 && y_pointer == 41)
||(x_pointer == 88 && y_pointer == 41)
||(x_pointer == 89 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 105 && y_pointer == 41)
||(x_pointer == 106 && y_pointer == 41)
||(x_pointer == 107 && y_pointer == 41)
||(x_pointer == 108 && y_pointer == 41)
||(x_pointer == 109 && y_pointer == 41)
||(x_pointer == 110 && y_pointer == 41)
||(x_pointer == 117 && y_pointer == 41)
||(x_pointer == 118 && y_pointer == 41)
||(x_pointer == 119 && y_pointer == 41)
||(x_pointer == 130 && y_pointer == 41)
||(x_pointer == 131 && y_pointer == 41)
||(x_pointer == 132 && y_pointer == 41)
||(x_pointer == 135 && y_pointer == 41)
||(x_pointer == 136 && y_pointer == 41)
||(x_pointer == 137 && y_pointer == 41)
||(x_pointer == 138 && y_pointer == 41)
||(x_pointer == 20 && y_pointer == 42)
||(x_pointer == 21 && y_pointer == 42)
||(x_pointer == 22 && y_pointer == 42)
||(x_pointer == 28 && y_pointer == 42)
||(x_pointer == 29 && y_pointer == 42)
||(x_pointer == 30 && y_pointer == 42)
||(x_pointer == 31 && y_pointer == 42)
||(x_pointer == 35 && y_pointer == 42)
||(x_pointer == 36 && y_pointer == 42)
||(x_pointer == 37 && y_pointer == 42)
||(x_pointer == 38 && y_pointer == 42)
||(x_pointer == 42 && y_pointer == 42)
||(x_pointer == 43 && y_pointer == 42)
||(x_pointer == 44 && y_pointer == 42)
||(x_pointer == 45 && y_pointer == 42)
||(x_pointer == 49 && y_pointer == 42)
||(x_pointer == 50 && y_pointer == 42)
||(x_pointer == 51 && y_pointer == 42)
||(x_pointer == 54 && y_pointer == 42)
||(x_pointer == 55 && y_pointer == 42)
||(x_pointer == 56 && y_pointer == 42)
||(x_pointer == 57 && y_pointer == 42)
||(x_pointer == 60 && y_pointer == 42)
||(x_pointer == 61 && y_pointer == 42)
||(x_pointer == 62 && y_pointer == 42)
||(x_pointer == 67 && y_pointer == 42)
||(x_pointer == 68 && y_pointer == 42)
||(x_pointer == 69 && y_pointer == 42)
||(x_pointer == 87 && y_pointer == 42)
||(x_pointer == 88 && y_pointer == 42)
||(x_pointer == 89 && y_pointer == 42)
||(x_pointer == 96 && y_pointer == 42)
||(x_pointer == 97 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 105 && y_pointer == 42)
||(x_pointer == 106 && y_pointer == 42)
||(x_pointer == 107 && y_pointer == 42)
||(x_pointer == 108 && y_pointer == 42)
||(x_pointer == 109 && y_pointer == 42)
||(x_pointer == 110 && y_pointer == 42)
||(x_pointer == 117 && y_pointer == 42)
||(x_pointer == 118 && y_pointer == 42)
||(x_pointer == 119 && y_pointer == 42)
||(x_pointer == 130 && y_pointer == 42)
||(x_pointer == 131 && y_pointer == 42)
||(x_pointer == 132 && y_pointer == 42)
||(x_pointer == 136 && y_pointer == 42)
||(x_pointer == 137 && y_pointer == 42)
||(x_pointer == 138 && y_pointer == 42)
||(x_pointer == 20 && y_pointer == 43)
||(x_pointer == 21 && y_pointer == 43)
||(x_pointer == 22 && y_pointer == 43)
||(x_pointer == 28 && y_pointer == 43)
||(x_pointer == 29 && y_pointer == 43)
||(x_pointer == 30 && y_pointer == 43)
||(x_pointer == 31 && y_pointer == 43)
||(x_pointer == 35 && y_pointer == 43)
||(x_pointer == 36 && y_pointer == 43)
||(x_pointer == 37 && y_pointer == 43)
||(x_pointer == 38 && y_pointer == 43)
||(x_pointer == 39 && y_pointer == 43)
||(x_pointer == 40 && y_pointer == 43)
||(x_pointer == 41 && y_pointer == 43)
||(x_pointer == 42 && y_pointer == 43)
||(x_pointer == 43 && y_pointer == 43)
||(x_pointer == 44 && y_pointer == 43)
||(x_pointer == 45 && y_pointer == 43)
||(x_pointer == 49 && y_pointer == 43)
||(x_pointer == 50 && y_pointer == 43)
||(x_pointer == 51 && y_pointer == 43)
||(x_pointer == 54 && y_pointer == 43)
||(x_pointer == 55 && y_pointer == 43)
||(x_pointer == 56 && y_pointer == 43)
||(x_pointer == 57 && y_pointer == 43)
||(x_pointer == 60 && y_pointer == 43)
||(x_pointer == 61 && y_pointer == 43)
||(x_pointer == 62 && y_pointer == 43)
||(x_pointer == 67 && y_pointer == 43)
||(x_pointer == 68 && y_pointer == 43)
||(x_pointer == 69 && y_pointer == 43)
||(x_pointer == 87 && y_pointer == 43)
||(x_pointer == 88 && y_pointer == 43)
||(x_pointer == 89 && y_pointer == 43)
||(x_pointer == 96 && y_pointer == 43)
||(x_pointer == 97 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 105 && y_pointer == 43)
||(x_pointer == 106 && y_pointer == 43)
||(x_pointer == 107 && y_pointer == 43)
||(x_pointer == 108 && y_pointer == 43)
||(x_pointer == 109 && y_pointer == 43)
||(x_pointer == 110 && y_pointer == 43)
||(x_pointer == 117 && y_pointer == 43)
||(x_pointer == 118 && y_pointer == 43)
||(x_pointer == 119 && y_pointer == 43)
||(x_pointer == 130 && y_pointer == 43)
||(x_pointer == 131 && y_pointer == 43)
||(x_pointer == 132 && y_pointer == 43)
||(x_pointer == 136 && y_pointer == 43)
||(x_pointer == 137 && y_pointer == 43)
||(x_pointer == 138 && y_pointer == 43)
||(x_pointer == 139 && y_pointer == 43)
||(x_pointer == 20 && y_pointer == 44)
||(x_pointer == 21 && y_pointer == 44)
||(x_pointer == 22 && y_pointer == 44)
||(x_pointer == 28 && y_pointer == 44)
||(x_pointer == 29 && y_pointer == 44)
||(x_pointer == 30 && y_pointer == 44)
||(x_pointer == 31 && y_pointer == 44)
||(x_pointer == 35 && y_pointer == 44)
||(x_pointer == 36 && y_pointer == 44)
||(x_pointer == 37 && y_pointer == 44)
||(x_pointer == 38 && y_pointer == 44)
||(x_pointer == 39 && y_pointer == 44)
||(x_pointer == 40 && y_pointer == 44)
||(x_pointer == 41 && y_pointer == 44)
||(x_pointer == 42 && y_pointer == 44)
||(x_pointer == 43 && y_pointer == 44)
||(x_pointer == 44 && y_pointer == 44)
||(x_pointer == 45 && y_pointer == 44)
||(x_pointer == 49 && y_pointer == 44)
||(x_pointer == 50 && y_pointer == 44)
||(x_pointer == 51 && y_pointer == 44)
||(x_pointer == 54 && y_pointer == 44)
||(x_pointer == 55 && y_pointer == 44)
||(x_pointer == 56 && y_pointer == 44)
||(x_pointer == 57 && y_pointer == 44)
||(x_pointer == 60 && y_pointer == 44)
||(x_pointer == 61 && y_pointer == 44)
||(x_pointer == 62 && y_pointer == 44)
||(x_pointer == 67 && y_pointer == 44)
||(x_pointer == 68 && y_pointer == 44)
||(x_pointer == 69 && y_pointer == 44)
||(x_pointer == 87 && y_pointer == 44)
||(x_pointer == 88 && y_pointer == 44)
||(x_pointer == 89 && y_pointer == 44)
||(x_pointer == 96 && y_pointer == 44)
||(x_pointer == 97 && y_pointer == 44)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 105 && y_pointer == 44)
||(x_pointer == 106 && y_pointer == 44)
||(x_pointer == 107 && y_pointer == 44)
||(x_pointer == 108 && y_pointer == 44)
||(x_pointer == 109 && y_pointer == 44)
||(x_pointer == 110 && y_pointer == 44)
||(x_pointer == 117 && y_pointer == 44)
||(x_pointer == 118 && y_pointer == 44)
||(x_pointer == 119 && y_pointer == 44)
||(x_pointer == 130 && y_pointer == 44)
||(x_pointer == 131 && y_pointer == 44)
||(x_pointer == 132 && y_pointer == 44)
||(x_pointer == 137 && y_pointer == 44)
||(x_pointer == 138 && y_pointer == 44)
||(x_pointer == 139 && y_pointer == 44)
||(x_pointer == 20 && y_pointer == 45)
||(x_pointer == 21 && y_pointer == 45)
||(x_pointer == 22 && y_pointer == 45)
||(x_pointer == 28 && y_pointer == 45)
||(x_pointer == 29 && y_pointer == 45)
||(x_pointer == 30 && y_pointer == 45)
||(x_pointer == 31 && y_pointer == 45)
||(x_pointer == 34 && y_pointer == 45)
||(x_pointer == 35 && y_pointer == 45)
||(x_pointer == 36 && y_pointer == 45)
||(x_pointer == 37 && y_pointer == 45)
||(x_pointer == 43 && y_pointer == 45)
||(x_pointer == 44 && y_pointer == 45)
||(x_pointer == 45 && y_pointer == 45)
||(x_pointer == 46 && y_pointer == 45)
||(x_pointer == 49 && y_pointer == 45)
||(x_pointer == 50 && y_pointer == 45)
||(x_pointer == 51 && y_pointer == 45)
||(x_pointer == 55 && y_pointer == 45)
||(x_pointer == 56 && y_pointer == 45)
||(x_pointer == 60 && y_pointer == 45)
||(x_pointer == 61 && y_pointer == 45)
||(x_pointer == 62 && y_pointer == 45)
||(x_pointer == 67 && y_pointer == 45)
||(x_pointer == 68 && y_pointer == 45)
||(x_pointer == 69 && y_pointer == 45)
||(x_pointer == 87 && y_pointer == 45)
||(x_pointer == 88 && y_pointer == 45)
||(x_pointer == 89 && y_pointer == 45)
||(x_pointer == 96 && y_pointer == 45)
||(x_pointer == 97 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 106 && y_pointer == 45)
||(x_pointer == 107 && y_pointer == 45)
||(x_pointer == 108 && y_pointer == 45)
||(x_pointer == 109 && y_pointer == 45)
||(x_pointer == 117 && y_pointer == 45)
||(x_pointer == 118 && y_pointer == 45)
||(x_pointer == 119 && y_pointer == 45)
||(x_pointer == 130 && y_pointer == 45)
||(x_pointer == 131 && y_pointer == 45)
||(x_pointer == 132 && y_pointer == 45)
||(x_pointer == 137 && y_pointer == 45)
||(x_pointer == 138 && y_pointer == 45)
||(x_pointer == 139 && y_pointer == 45)
||(x_pointer == 140 && y_pointer == 45)
||(x_pointer == 20 && y_pointer == 46)
||(x_pointer == 21 && y_pointer == 46)
||(x_pointer == 22 && y_pointer == 46)
||(x_pointer == 28 && y_pointer == 46)
||(x_pointer == 29 && y_pointer == 46)
||(x_pointer == 30 && y_pointer == 46)
||(x_pointer == 31 && y_pointer == 46)
||(x_pointer == 34 && y_pointer == 46)
||(x_pointer == 35 && y_pointer == 46)
||(x_pointer == 36 && y_pointer == 46)
||(x_pointer == 37 && y_pointer == 46)
||(x_pointer == 43 && y_pointer == 46)
||(x_pointer == 44 && y_pointer == 46)
||(x_pointer == 45 && y_pointer == 46)
||(x_pointer == 46 && y_pointer == 46)
||(x_pointer == 49 && y_pointer == 46)
||(x_pointer == 50 && y_pointer == 46)
||(x_pointer == 51 && y_pointer == 46)
||(x_pointer == 55 && y_pointer == 46)
||(x_pointer == 56 && y_pointer == 46)
||(x_pointer == 60 && y_pointer == 46)
||(x_pointer == 61 && y_pointer == 46)
||(x_pointer == 62 && y_pointer == 46)
||(x_pointer == 67 && y_pointer == 46)
||(x_pointer == 68 && y_pointer == 46)
||(x_pointer == 69 && y_pointer == 46)
||(x_pointer == 87 && y_pointer == 46)
||(x_pointer == 88 && y_pointer == 46)
||(x_pointer == 89 && y_pointer == 46)
||(x_pointer == 96 && y_pointer == 46)
||(x_pointer == 97 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 106 && y_pointer == 46)
||(x_pointer == 107 && y_pointer == 46)
||(x_pointer == 108 && y_pointer == 46)
||(x_pointer == 109 && y_pointer == 46)
||(x_pointer == 117 && y_pointer == 46)
||(x_pointer == 118 && y_pointer == 46)
||(x_pointer == 119 && y_pointer == 46)
||(x_pointer == 130 && y_pointer == 46)
||(x_pointer == 131 && y_pointer == 46)
||(x_pointer == 132 && y_pointer == 46)
||(x_pointer == 138 && y_pointer == 46)
||(x_pointer == 139 && y_pointer == 46)
||(x_pointer == 140 && y_pointer == 46)
||(x_pointer == 20 && y_pointer == 47)
||(x_pointer == 21 && y_pointer == 47)
||(x_pointer == 22 && y_pointer == 47)
||(x_pointer == 23 && y_pointer == 47)
||(x_pointer == 24 && y_pointer == 47)
||(x_pointer == 25 && y_pointer == 47)
||(x_pointer == 26 && y_pointer == 47)
||(x_pointer == 27 && y_pointer == 47)
||(x_pointer == 28 && y_pointer == 47)
||(x_pointer == 29 && y_pointer == 47)
||(x_pointer == 30 && y_pointer == 47)
||(x_pointer == 31 && y_pointer == 47)
||(x_pointer == 34 && y_pointer == 47)
||(x_pointer == 35 && y_pointer == 47)
||(x_pointer == 36 && y_pointer == 47)
||(x_pointer == 44 && y_pointer == 47)
||(x_pointer == 45 && y_pointer == 47)
||(x_pointer == 46 && y_pointer == 47)
||(x_pointer == 49 && y_pointer == 47)
||(x_pointer == 50 && y_pointer == 47)
||(x_pointer == 51 && y_pointer == 47)
||(x_pointer == 60 && y_pointer == 47)
||(x_pointer == 61 && y_pointer == 47)
||(x_pointer == 62 && y_pointer == 47)
||(x_pointer == 67 && y_pointer == 47)
||(x_pointer == 68 && y_pointer == 47)
||(x_pointer == 69 && y_pointer == 47)
||(x_pointer == 70 && y_pointer == 47)
||(x_pointer == 71 && y_pointer == 47)
||(x_pointer == 72 && y_pointer == 47)
||(x_pointer == 73 && y_pointer == 47)
||(x_pointer == 74 && y_pointer == 47)
||(x_pointer == 75 && y_pointer == 47)
||(x_pointer == 76 && y_pointer == 47)
||(x_pointer == 87 && y_pointer == 47)
||(x_pointer == 88 && y_pointer == 47)
||(x_pointer == 89 && y_pointer == 47)
||(x_pointer == 90 && y_pointer == 47)
||(x_pointer == 91 && y_pointer == 47)
||(x_pointer == 92 && y_pointer == 47)
||(x_pointer == 93 && y_pointer == 47)
||(x_pointer == 94 && y_pointer == 47)
||(x_pointer == 95 && y_pointer == 47)
||(x_pointer == 96 && y_pointer == 47)
||(x_pointer == 97 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 106 && y_pointer == 47)
||(x_pointer == 107 && y_pointer == 47)
||(x_pointer == 108 && y_pointer == 47)
||(x_pointer == 109 && y_pointer == 47)
||(x_pointer == 117 && y_pointer == 47)
||(x_pointer == 118 && y_pointer == 47)
||(x_pointer == 119 && y_pointer == 47)
||(x_pointer == 120 && y_pointer == 47)
||(x_pointer == 121 && y_pointer == 47)
||(x_pointer == 122 && y_pointer == 47)
||(x_pointer == 123 && y_pointer == 47)
||(x_pointer == 124 && y_pointer == 47)
||(x_pointer == 125 && y_pointer == 47)
||(x_pointer == 126 && y_pointer == 47)
||(x_pointer == 130 && y_pointer == 47)
||(x_pointer == 131 && y_pointer == 47)
||(x_pointer == 132 && y_pointer == 47)
||(x_pointer == 138 && y_pointer == 47)
||(x_pointer == 139 && y_pointer == 47)
||(x_pointer == 140 && y_pointer == 47)
||(x_pointer == 141 && y_pointer == 47)
||(x_pointer == 20 && y_pointer == 48)
||(x_pointer == 21 && y_pointer == 48)
||(x_pointer == 22 && y_pointer == 48)
||(x_pointer == 23 && y_pointer == 48)
||(x_pointer == 24 && y_pointer == 48)
||(x_pointer == 25 && y_pointer == 48)
||(x_pointer == 26 && y_pointer == 48)
||(x_pointer == 27 && y_pointer == 48)
||(x_pointer == 28 && y_pointer == 48)
||(x_pointer == 29 && y_pointer == 48)
||(x_pointer == 30 && y_pointer == 48)
||(x_pointer == 31 && y_pointer == 48)
||(x_pointer == 34 && y_pointer == 48)
||(x_pointer == 35 && y_pointer == 48)
||(x_pointer == 36 && y_pointer == 48)
||(x_pointer == 44 && y_pointer == 48)
||(x_pointer == 45 && y_pointer == 48)
||(x_pointer == 46 && y_pointer == 48)
||(x_pointer == 49 && y_pointer == 48)
||(x_pointer == 50 && y_pointer == 48)
||(x_pointer == 51 && y_pointer == 48)
||(x_pointer == 60 && y_pointer == 48)
||(x_pointer == 61 && y_pointer == 48)
||(x_pointer == 62 && y_pointer == 48)
||(x_pointer == 67 && y_pointer == 48)
||(x_pointer == 68 && y_pointer == 48)
||(x_pointer == 69 && y_pointer == 48)
||(x_pointer == 70 && y_pointer == 48)
||(x_pointer == 71 && y_pointer == 48)
||(x_pointer == 72 && y_pointer == 48)
||(x_pointer == 73 && y_pointer == 48)
||(x_pointer == 74 && y_pointer == 48)
||(x_pointer == 75 && y_pointer == 48)
||(x_pointer == 76 && y_pointer == 48)
||(x_pointer == 87 && y_pointer == 48)
||(x_pointer == 88 && y_pointer == 48)
||(x_pointer == 89 && y_pointer == 48)
||(x_pointer == 90 && y_pointer == 48)
||(x_pointer == 91 && y_pointer == 48)
||(x_pointer == 92 && y_pointer == 48)
||(x_pointer == 93 && y_pointer == 48)
||(x_pointer == 94 && y_pointer == 48)
||(x_pointer == 95 && y_pointer == 48)
||(x_pointer == 96 && y_pointer == 48)
||(x_pointer == 97 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 48)
||(x_pointer == 106 && y_pointer == 48)
||(x_pointer == 107 && y_pointer == 48)
||(x_pointer == 108 && y_pointer == 48)
||(x_pointer == 109 && y_pointer == 48)
||(x_pointer == 117 && y_pointer == 48)
||(x_pointer == 118 && y_pointer == 48)
||(x_pointer == 119 && y_pointer == 48)
||(x_pointer == 120 && y_pointer == 48)
||(x_pointer == 121 && y_pointer == 48)
||(x_pointer == 122 && y_pointer == 48)
||(x_pointer == 123 && y_pointer == 48)
||(x_pointer == 124 && y_pointer == 48)
||(x_pointer == 125 && y_pointer == 48)
||(x_pointer == 126 && y_pointer == 48)
||(x_pointer == 130 && y_pointer == 48)
||(x_pointer == 131 && y_pointer == 48)
||(x_pointer == 132 && y_pointer == 48)
||(x_pointer == 139 && y_pointer == 48)
||(x_pointer == 140 && y_pointer == 48)
||(x_pointer == 141 && y_pointer == 48)
||(x_pointer == 30 && y_pointer == 64)
||(x_pointer == 31 && y_pointer == 64)
||(x_pointer == 32 && y_pointer == 64)
||(x_pointer == 36 && y_pointer == 64)
||(x_pointer == 37 && y_pointer == 64)
||(x_pointer == 38 && y_pointer == 64)
||(x_pointer == 30 && y_pointer == 65)
||(x_pointer == 31 && y_pointer == 65)
||(x_pointer == 32 && y_pointer == 65)
||(x_pointer == 36 && y_pointer == 65)
||(x_pointer == 37 && y_pointer == 65)
||(x_pointer == 38 && y_pointer == 65)
||(x_pointer == 30 && y_pointer == 66)
||(x_pointer == 31 && y_pointer == 66)
||(x_pointer == 32 && y_pointer == 66)
||(x_pointer == 36 && y_pointer == 66)
||(x_pointer == 37 && y_pointer == 66)
||(x_pointer == 38 && y_pointer == 66)
||(x_pointer == 59 && y_pointer == 66)
||(x_pointer == 60 && y_pointer == 66)
||(x_pointer == 61 && y_pointer == 66)
||(x_pointer == 62 && y_pointer == 66)
||(x_pointer == 63 && y_pointer == 66)
||(x_pointer == 64 && y_pointer == 66)
||(x_pointer == 31 && y_pointer == 67)
||(x_pointer == 32 && y_pointer == 67)
||(x_pointer == 33 && y_pointer == 67)
||(x_pointer == 35 && y_pointer == 67)
||(x_pointer == 36 && y_pointer == 67)
||(x_pointer == 37 && y_pointer == 67)
||(x_pointer == 59 && y_pointer == 67)
||(x_pointer == 60 && y_pointer == 67)
||(x_pointer == 63 && y_pointer == 67)
||(x_pointer == 64 && y_pointer == 67)
||(x_pointer == 32 && y_pointer == 68)
||(x_pointer == 33 && y_pointer == 68)
||(x_pointer == 35 && y_pointer == 68)
||(x_pointer == 36 && y_pointer == 68)
||(x_pointer == 59 && y_pointer == 68)
||(x_pointer == 60 && y_pointer == 68)
||(x_pointer == 61 && y_pointer == 68)
||(x_pointer == 63 && y_pointer == 68)
||(x_pointer == 64 && y_pointer == 68)
||(x_pointer == 32 && y_pointer == 69)
||(x_pointer == 33 && y_pointer == 69)
||(x_pointer == 34 && y_pointer == 69)
||(x_pointer == 35 && y_pointer == 69)
||(x_pointer == 36 && y_pointer == 69)
||(x_pointer == 60 && y_pointer == 69)
||(x_pointer == 61 && y_pointer == 69)
||(x_pointer == 62 && y_pointer == 69)
||(x_pointer == 33 && y_pointer == 70)
||(x_pointer == 34 && y_pointer == 70)
||(x_pointer == 35 && y_pointer == 70)
||(x_pointer == 38 && y_pointer == 70)
||(x_pointer == 39 && y_pointer == 70)
||(x_pointer == 40 && y_pointer == 70)
||(x_pointer == 41 && y_pointer == 70)
||(x_pointer == 42 && y_pointer == 70)
||(x_pointer == 44 && y_pointer == 70)
||(x_pointer == 45 && y_pointer == 70)
||(x_pointer == 47 && y_pointer == 70)
||(x_pointer == 48 && y_pointer == 70)
||(x_pointer == 50 && y_pointer == 70)
||(x_pointer == 51 && y_pointer == 70)
||(x_pointer == 52 && y_pointer == 70)
||(x_pointer == 53 && y_pointer == 70)
||(x_pointer == 54 && y_pointer == 70)
||(x_pointer == 61 && y_pointer == 70)
||(x_pointer == 62 && y_pointer == 70)
||(x_pointer == 63 && y_pointer == 70)
||(x_pointer == 66 && y_pointer == 70)
||(x_pointer == 67 && y_pointer == 70)
||(x_pointer == 68 && y_pointer == 70)
||(x_pointer == 69 && y_pointer == 70)
||(x_pointer == 70 && y_pointer == 70)
||(x_pointer == 72 && y_pointer == 70)
||(x_pointer == 73 && y_pointer == 70)
||(x_pointer == 74 && y_pointer == 70)
||(x_pointer == 75 && y_pointer == 70)
||(x_pointer == 76 && y_pointer == 70)
||(x_pointer == 78 && y_pointer == 70)
||(x_pointer == 79 && y_pointer == 70)
||(x_pointer == 80 && y_pointer == 70)
||(x_pointer == 81 && y_pointer == 70)
||(x_pointer == 82 && y_pointer == 70)
||(x_pointer == 84 && y_pointer == 70)
||(x_pointer == 85 && y_pointer == 70)
||(x_pointer == 86 && y_pointer == 70)
||(x_pointer == 87 && y_pointer == 70)
||(x_pointer == 88 && y_pointer == 70)
||(x_pointer == 33 && y_pointer == 71)
||(x_pointer == 34 && y_pointer == 71)
||(x_pointer == 35 && y_pointer == 71)
||(x_pointer == 38 && y_pointer == 71)
||(x_pointer == 39 && y_pointer == 71)
||(x_pointer == 41 && y_pointer == 71)
||(x_pointer == 42 && y_pointer == 71)
||(x_pointer == 44 && y_pointer == 71)
||(x_pointer == 45 && y_pointer == 71)
||(x_pointer == 47 && y_pointer == 71)
||(x_pointer == 48 && y_pointer == 71)
||(x_pointer == 50 && y_pointer == 71)
||(x_pointer == 51 && y_pointer == 71)
||(x_pointer == 52 && y_pointer == 71)
||(x_pointer == 53 && y_pointer == 71)
||(x_pointer == 54 && y_pointer == 71)
||(x_pointer == 62 && y_pointer == 71)
||(x_pointer == 63 && y_pointer == 71)
||(x_pointer == 64 && y_pointer == 71)
||(x_pointer == 66 && y_pointer == 71)
||(x_pointer == 67 && y_pointer == 71)
||(x_pointer == 69 && y_pointer == 71)
||(x_pointer == 70 && y_pointer == 71)
||(x_pointer == 72 && y_pointer == 71)
||(x_pointer == 73 && y_pointer == 71)
||(x_pointer == 75 && y_pointer == 71)
||(x_pointer == 76 && y_pointer == 71)
||(x_pointer == 78 && y_pointer == 71)
||(x_pointer == 79 && y_pointer == 71)
||(x_pointer == 80 && y_pointer == 71)
||(x_pointer == 81 && y_pointer == 71)
||(x_pointer == 82 && y_pointer == 71)
||(x_pointer == 84 && y_pointer == 71)
||(x_pointer == 85 && y_pointer == 71)
||(x_pointer == 87 && y_pointer == 71)
||(x_pointer == 88 && y_pointer == 71)
||(x_pointer == 90 && y_pointer == 71)
||(x_pointer == 91 && y_pointer == 71)
||(x_pointer == 33 && y_pointer == 72)
||(x_pointer == 34 && y_pointer == 72)
||(x_pointer == 35 && y_pointer == 72)
||(x_pointer == 38 && y_pointer == 72)
||(x_pointer == 39 && y_pointer == 72)
||(x_pointer == 41 && y_pointer == 72)
||(x_pointer == 42 && y_pointer == 72)
||(x_pointer == 44 && y_pointer == 72)
||(x_pointer == 45 && y_pointer == 72)
||(x_pointer == 47 && y_pointer == 72)
||(x_pointer == 48 && y_pointer == 72)
||(x_pointer == 50 && y_pointer == 72)
||(x_pointer == 51 && y_pointer == 72)
||(x_pointer == 63 && y_pointer == 72)
||(x_pointer == 64 && y_pointer == 72)
||(x_pointer == 66 && y_pointer == 72)
||(x_pointer == 67 && y_pointer == 72)
||(x_pointer == 72 && y_pointer == 72)
||(x_pointer == 73 && y_pointer == 72)
||(x_pointer == 75 && y_pointer == 72)
||(x_pointer == 76 && y_pointer == 72)
||(x_pointer == 78 && y_pointer == 72)
||(x_pointer == 79 && y_pointer == 72)
||(x_pointer == 84 && y_pointer == 72)
||(x_pointer == 85 && y_pointer == 72)
||(x_pointer == 86 && y_pointer == 72)
||(x_pointer == 87 && y_pointer == 72)
||(x_pointer == 88 && y_pointer == 72)
||(x_pointer == 33 && y_pointer == 73)
||(x_pointer == 34 && y_pointer == 73)
||(x_pointer == 35 && y_pointer == 73)
||(x_pointer == 38 && y_pointer == 73)
||(x_pointer == 39 && y_pointer == 73)
||(x_pointer == 41 && y_pointer == 73)
||(x_pointer == 42 && y_pointer == 73)
||(x_pointer == 44 && y_pointer == 73)
||(x_pointer == 45 && y_pointer == 73)
||(x_pointer == 47 && y_pointer == 73)
||(x_pointer == 48 && y_pointer == 73)
||(x_pointer == 50 && y_pointer == 73)
||(x_pointer == 51 && y_pointer == 73)
||(x_pointer == 59 && y_pointer == 73)
||(x_pointer == 60 && y_pointer == 73)
||(x_pointer == 63 && y_pointer == 73)
||(x_pointer == 64 && y_pointer == 73)
||(x_pointer == 66 && y_pointer == 73)
||(x_pointer == 67 && y_pointer == 73)
||(x_pointer == 72 && y_pointer == 73)
||(x_pointer == 73 && y_pointer == 73)
||(x_pointer == 75 && y_pointer == 73)
||(x_pointer == 76 && y_pointer == 73)
||(x_pointer == 78 && y_pointer == 73)
||(x_pointer == 79 && y_pointer == 73)
||(x_pointer == 84 && y_pointer == 73)
||(x_pointer == 85 && y_pointer == 73)
||(x_pointer == 33 && y_pointer == 74)
||(x_pointer == 34 && y_pointer == 74)
||(x_pointer == 35 && y_pointer == 74)
||(x_pointer == 38 && y_pointer == 74)
||(x_pointer == 39 && y_pointer == 74)
||(x_pointer == 41 && y_pointer == 74)
||(x_pointer == 42 && y_pointer == 74)
||(x_pointer == 44 && y_pointer == 74)
||(x_pointer == 45 && y_pointer == 74)
||(x_pointer == 47 && y_pointer == 74)
||(x_pointer == 48 && y_pointer == 74)
||(x_pointer == 50 && y_pointer == 74)
||(x_pointer == 51 && y_pointer == 74)
||(x_pointer == 59 && y_pointer == 74)
||(x_pointer == 60 && y_pointer == 74)
||(x_pointer == 63 && y_pointer == 74)
||(x_pointer == 64 && y_pointer == 74)
||(x_pointer == 66 && y_pointer == 74)
||(x_pointer == 67 && y_pointer == 74)
||(x_pointer == 69 && y_pointer == 74)
||(x_pointer == 70 && y_pointer == 74)
||(x_pointer == 72 && y_pointer == 74)
||(x_pointer == 73 && y_pointer == 74)
||(x_pointer == 75 && y_pointer == 74)
||(x_pointer == 76 && y_pointer == 74)
||(x_pointer == 78 && y_pointer == 74)
||(x_pointer == 79 && y_pointer == 74)
||(x_pointer == 84 && y_pointer == 74)
||(x_pointer == 85 && y_pointer == 74)
||(x_pointer == 87 && y_pointer == 74)
||(x_pointer == 88 && y_pointer == 74)
||(x_pointer == 33 && y_pointer == 75)
||(x_pointer == 34 && y_pointer == 75)
||(x_pointer == 35 && y_pointer == 75)
||(x_pointer == 38 && y_pointer == 75)
||(x_pointer == 39 && y_pointer == 75)
||(x_pointer == 40 && y_pointer == 75)
||(x_pointer == 41 && y_pointer == 75)
||(x_pointer == 42 && y_pointer == 75)
||(x_pointer == 44 && y_pointer == 75)
||(x_pointer == 45 && y_pointer == 75)
||(x_pointer == 46 && y_pointer == 75)
||(x_pointer == 47 && y_pointer == 75)
||(x_pointer == 48 && y_pointer == 75)
||(x_pointer == 50 && y_pointer == 75)
||(x_pointer == 51 && y_pointer == 75)
||(x_pointer == 59 && y_pointer == 75)
||(x_pointer == 60 && y_pointer == 75)
||(x_pointer == 61 && y_pointer == 75)
||(x_pointer == 62 && y_pointer == 75)
||(x_pointer == 63 && y_pointer == 75)
||(x_pointer == 64 && y_pointer == 75)
||(x_pointer == 66 && y_pointer == 75)
||(x_pointer == 67 && y_pointer == 75)
||(x_pointer == 68 && y_pointer == 75)
||(x_pointer == 69 && y_pointer == 75)
||(x_pointer == 70 && y_pointer == 75)
||(x_pointer == 72 && y_pointer == 75)
||(x_pointer == 73 && y_pointer == 75)
||(x_pointer == 74 && y_pointer == 75)
||(x_pointer == 75 && y_pointer == 75)
||(x_pointer == 76 && y_pointer == 75)
||(x_pointer == 78 && y_pointer == 75)
||(x_pointer == 79 && y_pointer == 75)
||(x_pointer == 84 && y_pointer == 75)
||(x_pointer == 85 && y_pointer == 75)
||(x_pointer == 86 && y_pointer == 75)
||(x_pointer == 87 && y_pointer == 75)
||(x_pointer == 88 && y_pointer == 75)
||(x_pointer == 90 && y_pointer == 75)
||(x_pointer == 91 && y_pointer == 75)
||(x_pointer == 34 && y_pointer == 81)
||(x_pointer == 35 && y_pointer == 81)
||(x_pointer == 38 && y_pointer == 81)
||(x_pointer == 39 && y_pointer == 81)
||(x_pointer == 50 && y_pointer == 81)
||(x_pointer == 51 && y_pointer == 81)
||(x_pointer == 59 && y_pointer == 81)
||(x_pointer == 60 && y_pointer == 81)
||(x_pointer == 61 && y_pointer == 81)
||(x_pointer == 62 && y_pointer == 81)
||(x_pointer == 63 && y_pointer == 81)
||(x_pointer == 64 && y_pointer == 81)
||(x_pointer == 34 && y_pointer == 82)
||(x_pointer == 35 && y_pointer == 82)
||(x_pointer == 38 && y_pointer == 82)
||(x_pointer == 39 && y_pointer == 82)
||(x_pointer == 41 && y_pointer == 82)
||(x_pointer == 42 && y_pointer == 82)
||(x_pointer == 50 && y_pointer == 82)
||(x_pointer == 51 && y_pointer == 82)
||(x_pointer == 59 && y_pointer == 82)
||(x_pointer == 60 && y_pointer == 82)
||(x_pointer == 63 && y_pointer == 82)
||(x_pointer == 64 && y_pointer == 82)
||(x_pointer == 34 && y_pointer == 83)
||(x_pointer == 35 && y_pointer == 83)
||(x_pointer == 38 && y_pointer == 83)
||(x_pointer == 39 && y_pointer == 83)
||(x_pointer == 41 && y_pointer == 83)
||(x_pointer == 42 && y_pointer == 83)
||(x_pointer == 50 && y_pointer == 83)
||(x_pointer == 51 && y_pointer == 83)
||(x_pointer == 59 && y_pointer == 83)
||(x_pointer == 60 && y_pointer == 83)
||(x_pointer == 61 && y_pointer == 83)
||(x_pointer == 63 && y_pointer == 83)
||(x_pointer == 64 && y_pointer == 83)
||(x_pointer == 34 && y_pointer == 84)
||(x_pointer == 35 && y_pointer == 84)
||(x_pointer == 38 && y_pointer == 84)
||(x_pointer == 39 && y_pointer == 84)
||(x_pointer == 50 && y_pointer == 84)
||(x_pointer == 51 && y_pointer == 84)
||(x_pointer == 60 && y_pointer == 84)
||(x_pointer == 61 && y_pointer == 84)
||(x_pointer == 62 && y_pointer == 84)
||(x_pointer == 34 && y_pointer == 85)
||(x_pointer == 35 && y_pointer == 85)
||(x_pointer == 36 && y_pointer == 85)
||(x_pointer == 37 && y_pointer == 85)
||(x_pointer == 38 && y_pointer == 85)
||(x_pointer == 39 && y_pointer == 85)
||(x_pointer == 41 && y_pointer == 85)
||(x_pointer == 42 && y_pointer == 85)
||(x_pointer == 44 && y_pointer == 85)
||(x_pointer == 45 && y_pointer == 85)
||(x_pointer == 46 && y_pointer == 85)
||(x_pointer == 47 && y_pointer == 85)
||(x_pointer == 48 && y_pointer == 85)
||(x_pointer == 50 && y_pointer == 85)
||(x_pointer == 51 && y_pointer == 85)
||(x_pointer == 52 && y_pointer == 85)
||(x_pointer == 53 && y_pointer == 85)
||(x_pointer == 54 && y_pointer == 85)
||(x_pointer == 61 && y_pointer == 85)
||(x_pointer == 62 && y_pointer == 85)
||(x_pointer == 63 && y_pointer == 85)
||(x_pointer == 66 && y_pointer == 85)
||(x_pointer == 67 && y_pointer == 85)
||(x_pointer == 68 && y_pointer == 85)
||(x_pointer == 69 && y_pointer == 85)
||(x_pointer == 70 && y_pointer == 85)
||(x_pointer == 72 && y_pointer == 85)
||(x_pointer == 73 && y_pointer == 85)
||(x_pointer == 74 && y_pointer == 85)
||(x_pointer == 75 && y_pointer == 85)
||(x_pointer == 76 && y_pointer == 85)
||(x_pointer == 78 && y_pointer == 85)
||(x_pointer == 79 && y_pointer == 85)
||(x_pointer == 80 && y_pointer == 85)
||(x_pointer == 81 && y_pointer == 85)
||(x_pointer == 82 && y_pointer == 85)
||(x_pointer == 84 && y_pointer == 85)
||(x_pointer == 85 && y_pointer == 85)
||(x_pointer == 86 && y_pointer == 85)
||(x_pointer == 87 && y_pointer == 85)
||(x_pointer == 88 && y_pointer == 85)
||(x_pointer == 34 && y_pointer == 86)
||(x_pointer == 35 && y_pointer == 86)
||(x_pointer == 38 && y_pointer == 86)
||(x_pointer == 39 && y_pointer == 86)
||(x_pointer == 41 && y_pointer == 86)
||(x_pointer == 42 && y_pointer == 86)
||(x_pointer == 44 && y_pointer == 86)
||(x_pointer == 45 && y_pointer == 86)
||(x_pointer == 47 && y_pointer == 86)
||(x_pointer == 48 && y_pointer == 86)
||(x_pointer == 50 && y_pointer == 86)
||(x_pointer == 51 && y_pointer == 86)
||(x_pointer == 52 && y_pointer == 86)
||(x_pointer == 53 && y_pointer == 86)
||(x_pointer == 54 && y_pointer == 86)
||(x_pointer == 62 && y_pointer == 86)
||(x_pointer == 63 && y_pointer == 86)
||(x_pointer == 64 && y_pointer == 86)
||(x_pointer == 66 && y_pointer == 86)
||(x_pointer == 67 && y_pointer == 86)
||(x_pointer == 69 && y_pointer == 86)
||(x_pointer == 70 && y_pointer == 86)
||(x_pointer == 72 && y_pointer == 86)
||(x_pointer == 73 && y_pointer == 86)
||(x_pointer == 75 && y_pointer == 86)
||(x_pointer == 76 && y_pointer == 86)
||(x_pointer == 78 && y_pointer == 86)
||(x_pointer == 79 && y_pointer == 86)
||(x_pointer == 80 && y_pointer == 86)
||(x_pointer == 81 && y_pointer == 86)
||(x_pointer == 82 && y_pointer == 86)
||(x_pointer == 84 && y_pointer == 86)
||(x_pointer == 85 && y_pointer == 86)
||(x_pointer == 87 && y_pointer == 86)
||(x_pointer == 88 && y_pointer == 86)
||(x_pointer == 90 && y_pointer == 86)
||(x_pointer == 91 && y_pointer == 86)
||(x_pointer == 34 && y_pointer == 87)
||(x_pointer == 35 && y_pointer == 87)
||(x_pointer == 38 && y_pointer == 87)
||(x_pointer == 39 && y_pointer == 87)
||(x_pointer == 41 && y_pointer == 87)
||(x_pointer == 42 && y_pointer == 87)
||(x_pointer == 44 && y_pointer == 87)
||(x_pointer == 45 && y_pointer == 87)
||(x_pointer == 47 && y_pointer == 87)
||(x_pointer == 48 && y_pointer == 87)
||(x_pointer == 50 && y_pointer == 87)
||(x_pointer == 51 && y_pointer == 87)
||(x_pointer == 53 && y_pointer == 87)
||(x_pointer == 54 && y_pointer == 87)
||(x_pointer == 63 && y_pointer == 87)
||(x_pointer == 64 && y_pointer == 87)
||(x_pointer == 66 && y_pointer == 87)
||(x_pointer == 67 && y_pointer == 87)
||(x_pointer == 72 && y_pointer == 87)
||(x_pointer == 73 && y_pointer == 87)
||(x_pointer == 75 && y_pointer == 87)
||(x_pointer == 76 && y_pointer == 87)
||(x_pointer == 78 && y_pointer == 87)
||(x_pointer == 79 && y_pointer == 87)
||(x_pointer == 84 && y_pointer == 87)
||(x_pointer == 85 && y_pointer == 87)
||(x_pointer == 86 && y_pointer == 87)
||(x_pointer == 87 && y_pointer == 87)
||(x_pointer == 88 && y_pointer == 87)
||(x_pointer == 34 && y_pointer == 88)
||(x_pointer == 35 && y_pointer == 88)
||(x_pointer == 38 && y_pointer == 88)
||(x_pointer == 39 && y_pointer == 88)
||(x_pointer == 41 && y_pointer == 88)
||(x_pointer == 42 && y_pointer == 88)
||(x_pointer == 44 && y_pointer == 88)
||(x_pointer == 45 && y_pointer == 88)
||(x_pointer == 47 && y_pointer == 88)
||(x_pointer == 48 && y_pointer == 88)
||(x_pointer == 50 && y_pointer == 88)
||(x_pointer == 51 && y_pointer == 88)
||(x_pointer == 53 && y_pointer == 88)
||(x_pointer == 54 && y_pointer == 88)
||(x_pointer == 59 && y_pointer == 88)
||(x_pointer == 60 && y_pointer == 88)
||(x_pointer == 61 && y_pointer == 88)
||(x_pointer == 63 && y_pointer == 88)
||(x_pointer == 64 && y_pointer == 88)
||(x_pointer == 66 && y_pointer == 88)
||(x_pointer == 67 && y_pointer == 88)
||(x_pointer == 72 && y_pointer == 88)
||(x_pointer == 73 && y_pointer == 88)
||(x_pointer == 75 && y_pointer == 88)
||(x_pointer == 76 && y_pointer == 88)
||(x_pointer == 78 && y_pointer == 88)
||(x_pointer == 79 && y_pointer == 88)
||(x_pointer == 84 && y_pointer == 88)
||(x_pointer == 85 && y_pointer == 88)
||(x_pointer == 34 && y_pointer == 89)
||(x_pointer == 35 && y_pointer == 89)
||(x_pointer == 38 && y_pointer == 89)
||(x_pointer == 39 && y_pointer == 89)
||(x_pointer == 41 && y_pointer == 89)
||(x_pointer == 42 && y_pointer == 89)
||(x_pointer == 44 && y_pointer == 89)
||(x_pointer == 45 && y_pointer == 89)
||(x_pointer == 47 && y_pointer == 89)
||(x_pointer == 48 && y_pointer == 89)
||(x_pointer == 50 && y_pointer == 89)
||(x_pointer == 51 && y_pointer == 89)
||(x_pointer == 53 && y_pointer == 89)
||(x_pointer == 54 && y_pointer == 89)
||(x_pointer == 59 && y_pointer == 89)
||(x_pointer == 60 && y_pointer == 89)
||(x_pointer == 61 && y_pointer == 89)
||(x_pointer == 63 && y_pointer == 89)
||(x_pointer == 64 && y_pointer == 89)
||(x_pointer == 66 && y_pointer == 89)
||(x_pointer == 67 && y_pointer == 89)
||(x_pointer == 69 && y_pointer == 89)
||(x_pointer == 70 && y_pointer == 89)
||(x_pointer == 72 && y_pointer == 89)
||(x_pointer == 73 && y_pointer == 89)
||(x_pointer == 75 && y_pointer == 89)
||(x_pointer == 76 && y_pointer == 89)
||(x_pointer == 78 && y_pointer == 89)
||(x_pointer == 79 && y_pointer == 89)
||(x_pointer == 84 && y_pointer == 89)
||(x_pointer == 85 && y_pointer == 89)
||(x_pointer == 87 && y_pointer == 89)
||(x_pointer == 88 && y_pointer == 89)
||(x_pointer == 34 && y_pointer == 90)
||(x_pointer == 35 && y_pointer == 90)
||(x_pointer == 38 && y_pointer == 90)
||(x_pointer == 39 && y_pointer == 90)
||(x_pointer == 41 && y_pointer == 90)
||(x_pointer == 42 && y_pointer == 90)
||(x_pointer == 44 && y_pointer == 90)
||(x_pointer == 45 && y_pointer == 90)
||(x_pointer == 46 && y_pointer == 90)
||(x_pointer == 47 && y_pointer == 90)
||(x_pointer == 48 && y_pointer == 90)
||(x_pointer == 50 && y_pointer == 90)
||(x_pointer == 51 && y_pointer == 90)
||(x_pointer == 53 && y_pointer == 90)
||(x_pointer == 54 && y_pointer == 90)
||(x_pointer == 59 && y_pointer == 90)
||(x_pointer == 60 && y_pointer == 90)
||(x_pointer == 61 && y_pointer == 90)
||(x_pointer == 62 && y_pointer == 90)
||(x_pointer == 63 && y_pointer == 90)
||(x_pointer == 64 && y_pointer == 90)
||(x_pointer == 66 && y_pointer == 90)
||(x_pointer == 67 && y_pointer == 90)
||(x_pointer == 68 && y_pointer == 90)
||(x_pointer == 69 && y_pointer == 90)
||(x_pointer == 70 && y_pointer == 90)
||(x_pointer == 72 && y_pointer == 90)
||(x_pointer == 73 && y_pointer == 90)
||(x_pointer == 74 && y_pointer == 90)
||(x_pointer == 75 && y_pointer == 90)
||(x_pointer == 76 && y_pointer == 90)
||(x_pointer == 78 && y_pointer == 90)
||(x_pointer == 79 && y_pointer == 90)
||(x_pointer == 84 && y_pointer == 90)
||(x_pointer == 85 && y_pointer == 90)
||(x_pointer == 86 && y_pointer == 90)
||(x_pointer == 87 && y_pointer == 90)
||(x_pointer == 88 && y_pointer == 90)
||(x_pointer == 90 && y_pointer == 90)
||(x_pointer == 91 && y_pointer == 90)
||(x_pointer == 47 && y_pointer == 91)
||(x_pointer == 48 && y_pointer == 91)
||(x_pointer == 44 && y_pointer == 92)
||(x_pointer == 45 && y_pointer == 92)
||(x_pointer == 46 && y_pointer == 92)
||(x_pointer == 47 && y_pointer == 92)
||(x_pointer == 48 && y_pointer == 92);
endmodule