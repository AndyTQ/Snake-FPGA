module game_barrier_setter(clk, ingame, current_level, x_pointer, y_pointer, barrier);
   input ingame;
	input [3:0] current_level;
   input clk;
   input [7:0]x_pointer;
	input [6:0]y_pointer;
	output reg barrier; 

	always@(posedge clk)
	begin
		if (ingame)
			 begin
			 if (barrier_pixel_0 || barrier_pixel_1 || barrier_pixel_2)
				 barrier <= 1'b1;
			 else
				 barrier <= 1'b0;
			 end
	end
	wire barrier_pixel_0 = 1'b0;
	wire barrier_pixel_1 = current_level == 1 && ((x_pointer == 30 && y_pointer == 60)
||(x_pointer == 31 && y_pointer == 60)
||(x_pointer == 32 && y_pointer == 60)
||(x_pointer == 33 && y_pointer == 60)
||(x_pointer == 34 && y_pointer == 60)
||(x_pointer == 35 && y_pointer == 60)
||(x_pointer == 36 && y_pointer == 60)
||(x_pointer == 37 && y_pointer == 60)
||(x_pointer == 38 && y_pointer == 60)
||(x_pointer == 39 && y_pointer == 60)
||(x_pointer == 40 && y_pointer == 60)
||(x_pointer == 41 && y_pointer == 60)
||(x_pointer == 42 && y_pointer == 60)
||(x_pointer == 43 && y_pointer == 60)
||(x_pointer == 44 && y_pointer == 60)
||(x_pointer == 45 && y_pointer == 60)
||(x_pointer == 46 && y_pointer == 60)
||(x_pointer == 47 && y_pointer == 60)
||(x_pointer == 48 && y_pointer == 60)
||(x_pointer == 49 && y_pointer == 60)
||(x_pointer == 50 && y_pointer == 60)
||(x_pointer == 51 && y_pointer == 60)
||(x_pointer == 52 && y_pointer == 60)
||(x_pointer == 53 && y_pointer == 60)
||(x_pointer == 54 && y_pointer == 60)
||(x_pointer == 55 && y_pointer == 60)
||(x_pointer == 56 && y_pointer == 60)
||(x_pointer == 57 && y_pointer == 60)
||(x_pointer == 58 && y_pointer == 60)
||(x_pointer == 59 && y_pointer == 60)
||(x_pointer == 60 && y_pointer == 60)
||(x_pointer == 61 && y_pointer == 60)
||(x_pointer == 62 && y_pointer == 60)
||(x_pointer == 97 && y_pointer == 60)
||(x_pointer == 98 && y_pointer == 60)
||(x_pointer == 99 && y_pointer == 60)
||(x_pointer == 100 && y_pointer == 60)
||(x_pointer == 101 && y_pointer == 60)
||(x_pointer == 102 && y_pointer == 60)
||(x_pointer == 103 && y_pointer == 60)
||(x_pointer == 104 && y_pointer == 60)
||(x_pointer == 105 && y_pointer == 60)
||(x_pointer == 106 && y_pointer == 60)
||(x_pointer == 107 && y_pointer == 60)
||(x_pointer == 108 && y_pointer == 60)
||(x_pointer == 109 && y_pointer == 60)
||(x_pointer == 110 && y_pointer == 60)
||(x_pointer == 111 && y_pointer == 60)
||(x_pointer == 112 && y_pointer == 60)
||(x_pointer == 113 && y_pointer == 60)
||(x_pointer == 114 && y_pointer == 60)
||(x_pointer == 115 && y_pointer == 60)
||(x_pointer == 116 && y_pointer == 60)
||(x_pointer == 117 && y_pointer == 60)
||(x_pointer == 118 && y_pointer == 60)
||(x_pointer == 119 && y_pointer == 60)
||(x_pointer == 120 && y_pointer == 60)
||(x_pointer == 121 && y_pointer == 60)
||(x_pointer == 122 && y_pointer == 60)
||(x_pointer == 123 && y_pointer == 60)
||(x_pointer == 124 && y_pointer == 60)
||(x_pointer == 125 && y_pointer == 60)
||(x_pointer == 126 && y_pointer == 60)
||(x_pointer == 127 && y_pointer == 60)
||(x_pointer == 128 && y_pointer == 60)
||(x_pointer == 129 && y_pointer == 60)
||(x_pointer == 30 && y_pointer == 61)
||(x_pointer == 31 && y_pointer == 61)
||(x_pointer == 32 && y_pointer == 61)
||(x_pointer == 33 && y_pointer == 61)
||(x_pointer == 34 && y_pointer == 61)
||(x_pointer == 35 && y_pointer == 61)
||(x_pointer == 36 && y_pointer == 61)
||(x_pointer == 37 && y_pointer == 61)
||(x_pointer == 38 && y_pointer == 61)
||(x_pointer == 39 && y_pointer == 61)
||(x_pointer == 40 && y_pointer == 61)
||(x_pointer == 41 && y_pointer == 61)
||(x_pointer == 42 && y_pointer == 61)
||(x_pointer == 43 && y_pointer == 61)
||(x_pointer == 44 && y_pointer == 61)
||(x_pointer == 45 && y_pointer == 61)
||(x_pointer == 46 && y_pointer == 61)
||(x_pointer == 47 && y_pointer == 61)
||(x_pointer == 48 && y_pointer == 61)
||(x_pointer == 49 && y_pointer == 61)
||(x_pointer == 50 && y_pointer == 61)
||(x_pointer == 51 && y_pointer == 61)
||(x_pointer == 52 && y_pointer == 61)
||(x_pointer == 53 && y_pointer == 61)
||(x_pointer == 54 && y_pointer == 61)
||(x_pointer == 55 && y_pointer == 61)
||(x_pointer == 56 && y_pointer == 61)
||(x_pointer == 57 && y_pointer == 61)
||(x_pointer == 58 && y_pointer == 61)
||(x_pointer == 59 && y_pointer == 61)
||(x_pointer == 60 && y_pointer == 61)
||(x_pointer == 61 && y_pointer == 61)
||(x_pointer == 62 && y_pointer == 61)
||(x_pointer == 97 && y_pointer == 61)
||(x_pointer == 98 && y_pointer == 61)
||(x_pointer == 99 && y_pointer == 61)
||(x_pointer == 100 && y_pointer == 61)
||(x_pointer == 101 && y_pointer == 61)
||(x_pointer == 102 && y_pointer == 61)
||(x_pointer == 103 && y_pointer == 61)
||(x_pointer == 104 && y_pointer == 61)
||(x_pointer == 105 && y_pointer == 61)
||(x_pointer == 106 && y_pointer == 61)
||(x_pointer == 107 && y_pointer == 61)
||(x_pointer == 108 && y_pointer == 61)
||(x_pointer == 109 && y_pointer == 61)
||(x_pointer == 110 && y_pointer == 61)
||(x_pointer == 111 && y_pointer == 61)
||(x_pointer == 112 && y_pointer == 61)
||(x_pointer == 113 && y_pointer == 61)
||(x_pointer == 114 && y_pointer == 61)
||(x_pointer == 115 && y_pointer == 61)
||(x_pointer == 116 && y_pointer == 61)
||(x_pointer == 117 && y_pointer == 61)
||(x_pointer == 118 && y_pointer == 61)
||(x_pointer == 119 && y_pointer == 61)
||(x_pointer == 120 && y_pointer == 61)
||(x_pointer == 121 && y_pointer == 61)
||(x_pointer == 122 && y_pointer == 61)
||(x_pointer == 123 && y_pointer == 61)
||(x_pointer == 124 && y_pointer == 61)
||(x_pointer == 125 && y_pointer == 61)
||(x_pointer == 126 && y_pointer == 61)
||(x_pointer == 127 && y_pointer == 61)
||(x_pointer == 128 && y_pointer == 61)
||(x_pointer == 129 && y_pointer == 61)
||(x_pointer == 30 && y_pointer == 62)
||(x_pointer == 31 && y_pointer == 62)
||(x_pointer == 32 && y_pointer == 62)
||(x_pointer == 33 && y_pointer == 62)
||(x_pointer == 34 && y_pointer == 62)
||(x_pointer == 35 && y_pointer == 62)
||(x_pointer == 36 && y_pointer == 62)
||(x_pointer == 37 && y_pointer == 62)
||(x_pointer == 38 && y_pointer == 62)
||(x_pointer == 39 && y_pointer == 62)
||(x_pointer == 40 && y_pointer == 62)
||(x_pointer == 41 && y_pointer == 62)
||(x_pointer == 42 && y_pointer == 62)
||(x_pointer == 43 && y_pointer == 62)
||(x_pointer == 44 && y_pointer == 62)
||(x_pointer == 45 && y_pointer == 62)
||(x_pointer == 46 && y_pointer == 62)
||(x_pointer == 47 && y_pointer == 62)
||(x_pointer == 48 && y_pointer == 62)
||(x_pointer == 49 && y_pointer == 62)
||(x_pointer == 50 && y_pointer == 62)
||(x_pointer == 51 && y_pointer == 62)
||(x_pointer == 52 && y_pointer == 62)
||(x_pointer == 53 && y_pointer == 62)
||(x_pointer == 54 && y_pointer == 62)
||(x_pointer == 55 && y_pointer == 62)
||(x_pointer == 56 && y_pointer == 62)
||(x_pointer == 57 && y_pointer == 62)
||(x_pointer == 58 && y_pointer == 62)
||(x_pointer == 59 && y_pointer == 62)
||(x_pointer == 60 && y_pointer == 62)
||(x_pointer == 61 && y_pointer == 62)
||(x_pointer == 62 && y_pointer == 62)
||(x_pointer == 97 && y_pointer == 62)
||(x_pointer == 98 && y_pointer == 62)
||(x_pointer == 99 && y_pointer == 62)
||(x_pointer == 100 && y_pointer == 62)
||(x_pointer == 101 && y_pointer == 62)
||(x_pointer == 102 && y_pointer == 62)
||(x_pointer == 103 && y_pointer == 62)
||(x_pointer == 104 && y_pointer == 62)
||(x_pointer == 105 && y_pointer == 62)
||(x_pointer == 106 && y_pointer == 62)
||(x_pointer == 107 && y_pointer == 62)
||(x_pointer == 108 && y_pointer == 62)
||(x_pointer == 109 && y_pointer == 62)
||(x_pointer == 110 && y_pointer == 62)
||(x_pointer == 111 && y_pointer == 62)
||(x_pointer == 112 && y_pointer == 62)
||(x_pointer == 113 && y_pointer == 62)
||(x_pointer == 114 && y_pointer == 62)
||(x_pointer == 115 && y_pointer == 62)
||(x_pointer == 116 && y_pointer == 62)
||(x_pointer == 117 && y_pointer == 62)
||(x_pointer == 118 && y_pointer == 62)
||(x_pointer == 119 && y_pointer == 62)
||(x_pointer == 120 && y_pointer == 62)
||(x_pointer == 121 && y_pointer == 62)
||(x_pointer == 122 && y_pointer == 62)
||(x_pointer == 123 && y_pointer == 62)
||(x_pointer == 124 && y_pointer == 62)
||(x_pointer == 125 && y_pointer == 62)
||(x_pointer == 126 && y_pointer == 62)
||(x_pointer == 127 && y_pointer == 62)
||(x_pointer == 128 && y_pointer == 62)
||(x_pointer == 129 && y_pointer == 62)
||(x_pointer == 30 && y_pointer == 63)
||(x_pointer == 31 && y_pointer == 63)
||(x_pointer == 32 && y_pointer == 63)
||(x_pointer == 33 && y_pointer == 63)
||(x_pointer == 34 && y_pointer == 63)
||(x_pointer == 35 && y_pointer == 63)
||(x_pointer == 36 && y_pointer == 63)
||(x_pointer == 37 && y_pointer == 63)
||(x_pointer == 38 && y_pointer == 63)
||(x_pointer == 39 && y_pointer == 63)
||(x_pointer == 40 && y_pointer == 63)
||(x_pointer == 41 && y_pointer == 63)
||(x_pointer == 42 && y_pointer == 63)
||(x_pointer == 43 && y_pointer == 63)
||(x_pointer == 44 && y_pointer == 63)
||(x_pointer == 45 && y_pointer == 63)
||(x_pointer == 46 && y_pointer == 63)
||(x_pointer == 47 && y_pointer == 63)
||(x_pointer == 48 && y_pointer == 63)
||(x_pointer == 49 && y_pointer == 63)
||(x_pointer == 50 && y_pointer == 63)
||(x_pointer == 51 && y_pointer == 63)
||(x_pointer == 52 && y_pointer == 63)
||(x_pointer == 53 && y_pointer == 63)
||(x_pointer == 54 && y_pointer == 63)
||(x_pointer == 55 && y_pointer == 63)
||(x_pointer == 56 && y_pointer == 63)
||(x_pointer == 57 && y_pointer == 63)
||(x_pointer == 58 && y_pointer == 63)
||(x_pointer == 59 && y_pointer == 63)
||(x_pointer == 60 && y_pointer == 63)
||(x_pointer == 61 && y_pointer == 63)
||(x_pointer == 62 && y_pointer == 63)
||(x_pointer == 97 && y_pointer == 63)
||(x_pointer == 98 && y_pointer == 63)
||(x_pointer == 99 && y_pointer == 63)
||(x_pointer == 100 && y_pointer == 63)
||(x_pointer == 101 && y_pointer == 63)
||(x_pointer == 102 && y_pointer == 63)
||(x_pointer == 103 && y_pointer == 63)
||(x_pointer == 104 && y_pointer == 63)
||(x_pointer == 105 && y_pointer == 63)
||(x_pointer == 106 && y_pointer == 63)
||(x_pointer == 107 && y_pointer == 63)
||(x_pointer == 108 && y_pointer == 63)
||(x_pointer == 109 && y_pointer == 63)
||(x_pointer == 110 && y_pointer == 63)
||(x_pointer == 111 && y_pointer == 63)
||(x_pointer == 112 && y_pointer == 63)
||(x_pointer == 113 && y_pointer == 63)
||(x_pointer == 114 && y_pointer == 63)
||(x_pointer == 115 && y_pointer == 63)
||(x_pointer == 116 && y_pointer == 63)
||(x_pointer == 117 && y_pointer == 63)
||(x_pointer == 118 && y_pointer == 63)
||(x_pointer == 119 && y_pointer == 63)
||(x_pointer == 120 && y_pointer == 63)
||(x_pointer == 121 && y_pointer == 63)
||(x_pointer == 122 && y_pointer == 63)
||(x_pointer == 123 && y_pointer == 63)
||(x_pointer == 124 && y_pointer == 63)
||(x_pointer == 125 && y_pointer == 63)
||(x_pointer == 126 && y_pointer == 63)
||(x_pointer == 127 && y_pointer == 63)
||(x_pointer == 128 && y_pointer == 63)
||(x_pointer == 129 && y_pointer == 63)
||(x_pointer == 30 && y_pointer == 64)
||(x_pointer == 31 && y_pointer == 64)
||(x_pointer == 32 && y_pointer == 64)
||(x_pointer == 33 && y_pointer == 64)
||(x_pointer == 34 && y_pointer == 64)
||(x_pointer == 35 && y_pointer == 64)
||(x_pointer == 36 && y_pointer == 64)
||(x_pointer == 37 && y_pointer == 64)
||(x_pointer == 38 && y_pointer == 64)
||(x_pointer == 39 && y_pointer == 64)
||(x_pointer == 40 && y_pointer == 64)
||(x_pointer == 41 && y_pointer == 64)
||(x_pointer == 42 && y_pointer == 64)
||(x_pointer == 43 && y_pointer == 64)
||(x_pointer == 44 && y_pointer == 64)
||(x_pointer == 45 && y_pointer == 64)
||(x_pointer == 46 && y_pointer == 64)
||(x_pointer == 47 && y_pointer == 64)
||(x_pointer == 48 && y_pointer == 64)
||(x_pointer == 49 && y_pointer == 64)
||(x_pointer == 50 && y_pointer == 64)
||(x_pointer == 51 && y_pointer == 64)
||(x_pointer == 52 && y_pointer == 64)
||(x_pointer == 53 && y_pointer == 64)
||(x_pointer == 54 && y_pointer == 64)
||(x_pointer == 55 && y_pointer == 64)
||(x_pointer == 56 && y_pointer == 64)
||(x_pointer == 57 && y_pointer == 64)
||(x_pointer == 58 && y_pointer == 64)
||(x_pointer == 59 && y_pointer == 64)
||(x_pointer == 60 && y_pointer == 64)
||(x_pointer == 61 && y_pointer == 64)
||(x_pointer == 62 && y_pointer == 64)
||(x_pointer == 97 && y_pointer == 64)
||(x_pointer == 98 && y_pointer == 64)
||(x_pointer == 99 && y_pointer == 64)
||(x_pointer == 100 && y_pointer == 64)
||(x_pointer == 101 && y_pointer == 64)
||(x_pointer == 102 && y_pointer == 64)
||(x_pointer == 103 && y_pointer == 64)
||(x_pointer == 104 && y_pointer == 64)
||(x_pointer == 105 && y_pointer == 64)
||(x_pointer == 106 && y_pointer == 64)
||(x_pointer == 107 && y_pointer == 64)
||(x_pointer == 108 && y_pointer == 64)
||(x_pointer == 109 && y_pointer == 64)
||(x_pointer == 110 && y_pointer == 64)
||(x_pointer == 111 && y_pointer == 64)
||(x_pointer == 112 && y_pointer == 64)
||(x_pointer == 113 && y_pointer == 64)
||(x_pointer == 114 && y_pointer == 64)
||(x_pointer == 115 && y_pointer == 64)
||(x_pointer == 116 && y_pointer == 64)
||(x_pointer == 117 && y_pointer == 64)
||(x_pointer == 118 && y_pointer == 64)
||(x_pointer == 119 && y_pointer == 64)
||(x_pointer == 120 && y_pointer == 64)
||(x_pointer == 121 && y_pointer == 64)
||(x_pointer == 122 && y_pointer == 64)
||(x_pointer == 123 && y_pointer == 64)
||(x_pointer == 124 && y_pointer == 64)
||(x_pointer == 125 && y_pointer == 64)
||(x_pointer == 126 && y_pointer == 64)
||(x_pointer == 127 && y_pointer == 64)
||(x_pointer == 128 && y_pointer == 64)
||(x_pointer == 129 && y_pointer == 64)
||(x_pointer == 30 && y_pointer == 65)
||(x_pointer == 31 && y_pointer == 65)
||(x_pointer == 32 && y_pointer == 65)
||(x_pointer == 33 && y_pointer == 65)
||(x_pointer == 34 && y_pointer == 65)
||(x_pointer == 35 && y_pointer == 65)
||(x_pointer == 36 && y_pointer == 65)
||(x_pointer == 37 && y_pointer == 65)
||(x_pointer == 38 && y_pointer == 65)
||(x_pointer == 39 && y_pointer == 65)
||(x_pointer == 40 && y_pointer == 65)
||(x_pointer == 41 && y_pointer == 65)
||(x_pointer == 42 && y_pointer == 65)
||(x_pointer == 43 && y_pointer == 65)
||(x_pointer == 44 && y_pointer == 65)
||(x_pointer == 45 && y_pointer == 65)
||(x_pointer == 46 && y_pointer == 65)
||(x_pointer == 47 && y_pointer == 65)
||(x_pointer == 48 && y_pointer == 65)
||(x_pointer == 49 && y_pointer == 65)
||(x_pointer == 50 && y_pointer == 65)
||(x_pointer == 51 && y_pointer == 65)
||(x_pointer == 52 && y_pointer == 65)
||(x_pointer == 53 && y_pointer == 65)
||(x_pointer == 54 && y_pointer == 65)
||(x_pointer == 55 && y_pointer == 65)
||(x_pointer == 56 && y_pointer == 65)
||(x_pointer == 57 && y_pointer == 65)
||(x_pointer == 58 && y_pointer == 65)
||(x_pointer == 59 && y_pointer == 65)
||(x_pointer == 60 && y_pointer == 65)
||(x_pointer == 61 && y_pointer == 65)
||(x_pointer == 62 && y_pointer == 65)
||(x_pointer == 97 && y_pointer == 65)
||(x_pointer == 98 && y_pointer == 65)
||(x_pointer == 99 && y_pointer == 65)
||(x_pointer == 100 && y_pointer == 65)
||(x_pointer == 101 && y_pointer == 65)
||(x_pointer == 102 && y_pointer == 65)
||(x_pointer == 103 && y_pointer == 65)
||(x_pointer == 104 && y_pointer == 65)
||(x_pointer == 105 && y_pointer == 65)
||(x_pointer == 106 && y_pointer == 65)
||(x_pointer == 107 && y_pointer == 65)
||(x_pointer == 108 && y_pointer == 65)
||(x_pointer == 109 && y_pointer == 65)
||(x_pointer == 110 && y_pointer == 65)
||(x_pointer == 111 && y_pointer == 65)
||(x_pointer == 112 && y_pointer == 65)
||(x_pointer == 113 && y_pointer == 65)
||(x_pointer == 114 && y_pointer == 65)
||(x_pointer == 115 && y_pointer == 65)
||(x_pointer == 116 && y_pointer == 65)
||(x_pointer == 117 && y_pointer == 65)
||(x_pointer == 118 && y_pointer == 65)
||(x_pointer == 119 && y_pointer == 65)
||(x_pointer == 120 && y_pointer == 65)
||(x_pointer == 121 && y_pointer == 65)
||(x_pointer == 122 && y_pointer == 65)
||(x_pointer == 123 && y_pointer == 65)
||(x_pointer == 124 && y_pointer == 65)
||(x_pointer == 125 && y_pointer == 65)
||(x_pointer == 126 && y_pointer == 65)
||(x_pointer == 127 && y_pointer == 65)
||(x_pointer == 128 && y_pointer == 65)
||(x_pointer == 129 && y_pointer == 65)
||(x_pointer == 30 && y_pointer == 66)
||(x_pointer == 31 && y_pointer == 66)
||(x_pointer == 32 && y_pointer == 66)
||(x_pointer == 33 && y_pointer == 66)
||(x_pointer == 34 && y_pointer == 66)
||(x_pointer == 35 && y_pointer == 66)
||(x_pointer == 36 && y_pointer == 66)
||(x_pointer == 37 && y_pointer == 66)
||(x_pointer == 38 && y_pointer == 66)
||(x_pointer == 39 && y_pointer == 66)
||(x_pointer == 40 && y_pointer == 66)
||(x_pointer == 41 && y_pointer == 66)
||(x_pointer == 42 && y_pointer == 66)
||(x_pointer == 43 && y_pointer == 66)
||(x_pointer == 44 && y_pointer == 66)
||(x_pointer == 45 && y_pointer == 66)
||(x_pointer == 46 && y_pointer == 66)
||(x_pointer == 47 && y_pointer == 66)
||(x_pointer == 48 && y_pointer == 66)
||(x_pointer == 49 && y_pointer == 66)
||(x_pointer == 50 && y_pointer == 66)
||(x_pointer == 51 && y_pointer == 66)
||(x_pointer == 52 && y_pointer == 66)
||(x_pointer == 53 && y_pointer == 66)
||(x_pointer == 54 && y_pointer == 66)
||(x_pointer == 55 && y_pointer == 66)
||(x_pointer == 56 && y_pointer == 66)
||(x_pointer == 57 && y_pointer == 66)
||(x_pointer == 58 && y_pointer == 66)
||(x_pointer == 59 && y_pointer == 66)
||(x_pointer == 60 && y_pointer == 66)
||(x_pointer == 61 && y_pointer == 66)
||(x_pointer == 62 && y_pointer == 66)
||(x_pointer == 97 && y_pointer == 66)
||(x_pointer == 98 && y_pointer == 66)
||(x_pointer == 99 && y_pointer == 66)
||(x_pointer == 100 && y_pointer == 66)
||(x_pointer == 101 && y_pointer == 66)
||(x_pointer == 102 && y_pointer == 66)
||(x_pointer == 103 && y_pointer == 66)
||(x_pointer == 104 && y_pointer == 66)
||(x_pointer == 105 && y_pointer == 66)
||(x_pointer == 106 && y_pointer == 66)
||(x_pointer == 107 && y_pointer == 66)
||(x_pointer == 108 && y_pointer == 66)
||(x_pointer == 109 && y_pointer == 66)
||(x_pointer == 110 && y_pointer == 66)
||(x_pointer == 111 && y_pointer == 66)
||(x_pointer == 112 && y_pointer == 66)
||(x_pointer == 113 && y_pointer == 66)
||(x_pointer == 114 && y_pointer == 66)
||(x_pointer == 115 && y_pointer == 66)
||(x_pointer == 116 && y_pointer == 66)
||(x_pointer == 117 && y_pointer == 66)
||(x_pointer == 118 && y_pointer == 66)
||(x_pointer == 119 && y_pointer == 66)
||(x_pointer == 120 && y_pointer == 66)
||(x_pointer == 121 && y_pointer == 66)
||(x_pointer == 122 && y_pointer == 66)
||(x_pointer == 123 && y_pointer == 66)
||(x_pointer == 124 && y_pointer == 66)
||(x_pointer == 125 && y_pointer == 66)
||(x_pointer == 126 && y_pointer == 66)
||(x_pointer == 127 && y_pointer == 66)
||(x_pointer == 128 && y_pointer == 66)
||(x_pointer == 129 && y_pointer == 66)
||(x_pointer == 30 && y_pointer == 67)
||(x_pointer == 31 && y_pointer == 67)
||(x_pointer == 32 && y_pointer == 67)
||(x_pointer == 33 && y_pointer == 67)
||(x_pointer == 34 && y_pointer == 67)
||(x_pointer == 35 && y_pointer == 67)
||(x_pointer == 36 && y_pointer == 67)
||(x_pointer == 37 && y_pointer == 67)
||(x_pointer == 38 && y_pointer == 67)
||(x_pointer == 39 && y_pointer == 67)
||(x_pointer == 40 && y_pointer == 67)
||(x_pointer == 41 && y_pointer == 67)
||(x_pointer == 42 && y_pointer == 67)
||(x_pointer == 43 && y_pointer == 67)
||(x_pointer == 44 && y_pointer == 67)
||(x_pointer == 45 && y_pointer == 67)
||(x_pointer == 46 && y_pointer == 67)
||(x_pointer == 47 && y_pointer == 67)
||(x_pointer == 48 && y_pointer == 67)
||(x_pointer == 49 && y_pointer == 67)
||(x_pointer == 50 && y_pointer == 67)
||(x_pointer == 51 && y_pointer == 67)
||(x_pointer == 52 && y_pointer == 67)
||(x_pointer == 53 && y_pointer == 67)
||(x_pointer == 54 && y_pointer == 67)
||(x_pointer == 55 && y_pointer == 67)
||(x_pointer == 56 && y_pointer == 67)
||(x_pointer == 57 && y_pointer == 67)
||(x_pointer == 58 && y_pointer == 67)
||(x_pointer == 59 && y_pointer == 67)
||(x_pointer == 60 && y_pointer == 67)
||(x_pointer == 61 && y_pointer == 67)
||(x_pointer == 62 && y_pointer == 67)
||(x_pointer == 97 && y_pointer == 67)
||(x_pointer == 98 && y_pointer == 67)
||(x_pointer == 99 && y_pointer == 67)
||(x_pointer == 100 && y_pointer == 67)
||(x_pointer == 101 && y_pointer == 67)
||(x_pointer == 102 && y_pointer == 67)
||(x_pointer == 103 && y_pointer == 67)
||(x_pointer == 104 && y_pointer == 67)
||(x_pointer == 105 && y_pointer == 67)
||(x_pointer == 106 && y_pointer == 67)
||(x_pointer == 107 && y_pointer == 67)
||(x_pointer == 108 && y_pointer == 67)
||(x_pointer == 109 && y_pointer == 67)
||(x_pointer == 110 && y_pointer == 67)
||(x_pointer == 111 && y_pointer == 67)
||(x_pointer == 112 && y_pointer == 67)
||(x_pointer == 113 && y_pointer == 67)
||(x_pointer == 114 && y_pointer == 67)
||(x_pointer == 115 && y_pointer == 67)
||(x_pointer == 116 && y_pointer == 67)
||(x_pointer == 117 && y_pointer == 67)
||(x_pointer == 118 && y_pointer == 67)
||(x_pointer == 119 && y_pointer == 67)
||(x_pointer == 120 && y_pointer == 67)
||(x_pointer == 121 && y_pointer == 67)
||(x_pointer == 122 && y_pointer == 67)
||(x_pointer == 123 && y_pointer == 67)
||(x_pointer == 124 && y_pointer == 67)
||(x_pointer == 125 && y_pointer == 67)
||(x_pointer == 126 && y_pointer == 67)
||(x_pointer == 127 && y_pointer == 67)
||(x_pointer == 128 && y_pointer == 67)
||(x_pointer == 129 && y_pointer == 67));
	wire barrier_pixel_2 = current_level == 2 && ((x_pointer == 43 && y_pointer == 21)
||(x_pointer == 44 && y_pointer == 21)
||(x_pointer == 45 && y_pointer == 21)
||(x_pointer == 46 && y_pointer == 21)
||(x_pointer == 47 && y_pointer == 21)
||(x_pointer == 48 && y_pointer == 21)
||(x_pointer == 49 && y_pointer == 21)
||(x_pointer == 50 && y_pointer == 21)
||(x_pointer == 51 && y_pointer == 21)
||(x_pointer == 52 && y_pointer == 21)
||(x_pointer == 53 && y_pointer == 21)
||(x_pointer == 54 && y_pointer == 21)
||(x_pointer == 55 && y_pointer == 21)
||(x_pointer == 56 && y_pointer == 21)
||(x_pointer == 57 && y_pointer == 21)
||(x_pointer == 58 && y_pointer == 21)
||(x_pointer == 59 && y_pointer == 21)
||(x_pointer == 60 && y_pointer == 21)
||(x_pointer == 61 && y_pointer == 21)
||(x_pointer == 62 && y_pointer == 21)
||(x_pointer == 63 && y_pointer == 21)
||(x_pointer == 64 && y_pointer == 21)
||(x_pointer == 65 && y_pointer == 21)
||(x_pointer == 66 && y_pointer == 21)
||(x_pointer == 67 && y_pointer == 21)
||(x_pointer == 68 && y_pointer == 21)
||(x_pointer == 69 && y_pointer == 21)
||(x_pointer == 70 && y_pointer == 21)
||(x_pointer == 90 && y_pointer == 21)
||(x_pointer == 91 && y_pointer == 21)
||(x_pointer == 92 && y_pointer == 21)
||(x_pointer == 93 && y_pointer == 21)
||(x_pointer == 94 && y_pointer == 21)
||(x_pointer == 95 && y_pointer == 21)
||(x_pointer == 96 && y_pointer == 21)
||(x_pointer == 97 && y_pointer == 21)
||(x_pointer == 98 && y_pointer == 21)
||(x_pointer == 99 && y_pointer == 21)
||(x_pointer == 100 && y_pointer == 21)
||(x_pointer == 101 && y_pointer == 21)
||(x_pointer == 102 && y_pointer == 21)
||(x_pointer == 103 && y_pointer == 21)
||(x_pointer == 104 && y_pointer == 21)
||(x_pointer == 105 && y_pointer == 21)
||(x_pointer == 106 && y_pointer == 21)
||(x_pointer == 107 && y_pointer == 21)
||(x_pointer == 108 && y_pointer == 21)
||(x_pointer == 109 && y_pointer == 21)
||(x_pointer == 110 && y_pointer == 21)
||(x_pointer == 111 && y_pointer == 21)
||(x_pointer == 112 && y_pointer == 21)
||(x_pointer == 113 && y_pointer == 21)
||(x_pointer == 114 && y_pointer == 21)
||(x_pointer == 115 && y_pointer == 21)
||(x_pointer == 116 && y_pointer == 21)
||(x_pointer == 117 && y_pointer == 21)
||(x_pointer == 43 && y_pointer == 22)
||(x_pointer == 44 && y_pointer == 22)
||(x_pointer == 45 && y_pointer == 22)
||(x_pointer == 46 && y_pointer == 22)
||(x_pointer == 47 && y_pointer == 22)
||(x_pointer == 48 && y_pointer == 22)
||(x_pointer == 49 && y_pointer == 22)
||(x_pointer == 50 && y_pointer == 22)
||(x_pointer == 51 && y_pointer == 22)
||(x_pointer == 52 && y_pointer == 22)
||(x_pointer == 53 && y_pointer == 22)
||(x_pointer == 54 && y_pointer == 22)
||(x_pointer == 55 && y_pointer == 22)
||(x_pointer == 56 && y_pointer == 22)
||(x_pointer == 57 && y_pointer == 22)
||(x_pointer == 58 && y_pointer == 22)
||(x_pointer == 59 && y_pointer == 22)
||(x_pointer == 60 && y_pointer == 22)
||(x_pointer == 61 && y_pointer == 22)
||(x_pointer == 62 && y_pointer == 22)
||(x_pointer == 63 && y_pointer == 22)
||(x_pointer == 64 && y_pointer == 22)
||(x_pointer == 65 && y_pointer == 22)
||(x_pointer == 66 && y_pointer == 22)
||(x_pointer == 67 && y_pointer == 22)
||(x_pointer == 68 && y_pointer == 22)
||(x_pointer == 69 && y_pointer == 22)
||(x_pointer == 70 && y_pointer == 22)
||(x_pointer == 90 && y_pointer == 22)
||(x_pointer == 91 && y_pointer == 22)
||(x_pointer == 92 && y_pointer == 22)
||(x_pointer == 93 && y_pointer == 22)
||(x_pointer == 94 && y_pointer == 22)
||(x_pointer == 95 && y_pointer == 22)
||(x_pointer == 96 && y_pointer == 22)
||(x_pointer == 97 && y_pointer == 22)
||(x_pointer == 98 && y_pointer == 22)
||(x_pointer == 99 && y_pointer == 22)
||(x_pointer == 100 && y_pointer == 22)
||(x_pointer == 101 && y_pointer == 22)
||(x_pointer == 102 && y_pointer == 22)
||(x_pointer == 103 && y_pointer == 22)
||(x_pointer == 104 && y_pointer == 22)
||(x_pointer == 105 && y_pointer == 22)
||(x_pointer == 106 && y_pointer == 22)
||(x_pointer == 107 && y_pointer == 22)
||(x_pointer == 108 && y_pointer == 22)
||(x_pointer == 109 && y_pointer == 22)
||(x_pointer == 110 && y_pointer == 22)
||(x_pointer == 111 && y_pointer == 22)
||(x_pointer == 112 && y_pointer == 22)
||(x_pointer == 113 && y_pointer == 22)
||(x_pointer == 114 && y_pointer == 22)
||(x_pointer == 115 && y_pointer == 22)
||(x_pointer == 116 && y_pointer == 22)
||(x_pointer == 117 && y_pointer == 22)
||(x_pointer == 43 && y_pointer == 23)
||(x_pointer == 44 && y_pointer == 23)
||(x_pointer == 45 && y_pointer == 23)
||(x_pointer == 46 && y_pointer == 23)
||(x_pointer == 47 && y_pointer == 23)
||(x_pointer == 48 && y_pointer == 23)
||(x_pointer == 49 && y_pointer == 23)
||(x_pointer == 50 && y_pointer == 23)
||(x_pointer == 51 && y_pointer == 23)
||(x_pointer == 52 && y_pointer == 23)
||(x_pointer == 53 && y_pointer == 23)
||(x_pointer == 54 && y_pointer == 23)
||(x_pointer == 55 && y_pointer == 23)
||(x_pointer == 56 && y_pointer == 23)
||(x_pointer == 57 && y_pointer == 23)
||(x_pointer == 58 && y_pointer == 23)
||(x_pointer == 59 && y_pointer == 23)
||(x_pointer == 60 && y_pointer == 23)
||(x_pointer == 61 && y_pointer == 23)
||(x_pointer == 62 && y_pointer == 23)
||(x_pointer == 63 && y_pointer == 23)
||(x_pointer == 64 && y_pointer == 23)
||(x_pointer == 65 && y_pointer == 23)
||(x_pointer == 66 && y_pointer == 23)
||(x_pointer == 67 && y_pointer == 23)
||(x_pointer == 68 && y_pointer == 23)
||(x_pointer == 69 && y_pointer == 23)
||(x_pointer == 70 && y_pointer == 23)
||(x_pointer == 90 && y_pointer == 23)
||(x_pointer == 91 && y_pointer == 23)
||(x_pointer == 92 && y_pointer == 23)
||(x_pointer == 93 && y_pointer == 23)
||(x_pointer == 94 && y_pointer == 23)
||(x_pointer == 95 && y_pointer == 23)
||(x_pointer == 96 && y_pointer == 23)
||(x_pointer == 97 && y_pointer == 23)
||(x_pointer == 98 && y_pointer == 23)
||(x_pointer == 99 && y_pointer == 23)
||(x_pointer == 100 && y_pointer == 23)
||(x_pointer == 101 && y_pointer == 23)
||(x_pointer == 102 && y_pointer == 23)
||(x_pointer == 103 && y_pointer == 23)
||(x_pointer == 104 && y_pointer == 23)
||(x_pointer == 105 && y_pointer == 23)
||(x_pointer == 106 && y_pointer == 23)
||(x_pointer == 107 && y_pointer == 23)
||(x_pointer == 108 && y_pointer == 23)
||(x_pointer == 109 && y_pointer == 23)
||(x_pointer == 110 && y_pointer == 23)
||(x_pointer == 111 && y_pointer == 23)
||(x_pointer == 112 && y_pointer == 23)
||(x_pointer == 113 && y_pointer == 23)
||(x_pointer == 114 && y_pointer == 23)
||(x_pointer == 115 && y_pointer == 23)
||(x_pointer == 116 && y_pointer == 23)
||(x_pointer == 117 && y_pointer == 23)
||(x_pointer == 43 && y_pointer == 24)
||(x_pointer == 44 && y_pointer == 24)
||(x_pointer == 45 && y_pointer == 24)
||(x_pointer == 46 && y_pointer == 24)
||(x_pointer == 47 && y_pointer == 24)
||(x_pointer == 48 && y_pointer == 24)
||(x_pointer == 49 && y_pointer == 24)
||(x_pointer == 50 && y_pointer == 24)
||(x_pointer == 51 && y_pointer == 24)
||(x_pointer == 52 && y_pointer == 24)
||(x_pointer == 53 && y_pointer == 24)
||(x_pointer == 54 && y_pointer == 24)
||(x_pointer == 55 && y_pointer == 24)
||(x_pointer == 56 && y_pointer == 24)
||(x_pointer == 57 && y_pointer == 24)
||(x_pointer == 58 && y_pointer == 24)
||(x_pointer == 59 && y_pointer == 24)
||(x_pointer == 60 && y_pointer == 24)
||(x_pointer == 61 && y_pointer == 24)
||(x_pointer == 62 && y_pointer == 24)
||(x_pointer == 63 && y_pointer == 24)
||(x_pointer == 64 && y_pointer == 24)
||(x_pointer == 65 && y_pointer == 24)
||(x_pointer == 66 && y_pointer == 24)
||(x_pointer == 67 && y_pointer == 24)
||(x_pointer == 68 && y_pointer == 24)
||(x_pointer == 69 && y_pointer == 24)
||(x_pointer == 70 && y_pointer == 24)
||(x_pointer == 90 && y_pointer == 24)
||(x_pointer == 91 && y_pointer == 24)
||(x_pointer == 92 && y_pointer == 24)
||(x_pointer == 93 && y_pointer == 24)
||(x_pointer == 94 && y_pointer == 24)
||(x_pointer == 95 && y_pointer == 24)
||(x_pointer == 96 && y_pointer == 24)
||(x_pointer == 97 && y_pointer == 24)
||(x_pointer == 98 && y_pointer == 24)
||(x_pointer == 99 && y_pointer == 24)
||(x_pointer == 100 && y_pointer == 24)
||(x_pointer == 101 && y_pointer == 24)
||(x_pointer == 102 && y_pointer == 24)
||(x_pointer == 103 && y_pointer == 24)
||(x_pointer == 104 && y_pointer == 24)
||(x_pointer == 105 && y_pointer == 24)
||(x_pointer == 106 && y_pointer == 24)
||(x_pointer == 107 && y_pointer == 24)
||(x_pointer == 108 && y_pointer == 24)
||(x_pointer == 109 && y_pointer == 24)
||(x_pointer == 110 && y_pointer == 24)
||(x_pointer == 111 && y_pointer == 24)
||(x_pointer == 112 && y_pointer == 24)
||(x_pointer == 113 && y_pointer == 24)
||(x_pointer == 114 && y_pointer == 24)
||(x_pointer == 115 && y_pointer == 24)
||(x_pointer == 116 && y_pointer == 24)
||(x_pointer == 117 && y_pointer == 24)
||(x_pointer == 43 && y_pointer == 25)
||(x_pointer == 44 && y_pointer == 25)
||(x_pointer == 45 && y_pointer == 25)
||(x_pointer == 46 && y_pointer == 25)
||(x_pointer == 47 && y_pointer == 25)
||(x_pointer == 48 && y_pointer == 25)
||(x_pointer == 49 && y_pointer == 25)
||(x_pointer == 50 && y_pointer == 25)
||(x_pointer == 51 && y_pointer == 25)
||(x_pointer == 52 && y_pointer == 25)
||(x_pointer == 53 && y_pointer == 25)
||(x_pointer == 54 && y_pointer == 25)
||(x_pointer == 55 && y_pointer == 25)
||(x_pointer == 56 && y_pointer == 25)
||(x_pointer == 57 && y_pointer == 25)
||(x_pointer == 58 && y_pointer == 25)
||(x_pointer == 59 && y_pointer == 25)
||(x_pointer == 60 && y_pointer == 25)
||(x_pointer == 61 && y_pointer == 25)
||(x_pointer == 62 && y_pointer == 25)
||(x_pointer == 63 && y_pointer == 25)
||(x_pointer == 64 && y_pointer == 25)
||(x_pointer == 65 && y_pointer == 25)
||(x_pointer == 66 && y_pointer == 25)
||(x_pointer == 67 && y_pointer == 25)
||(x_pointer == 68 && y_pointer == 25)
||(x_pointer == 69 && y_pointer == 25)
||(x_pointer == 70 && y_pointer == 25)
||(x_pointer == 90 && y_pointer == 25)
||(x_pointer == 91 && y_pointer == 25)
||(x_pointer == 92 && y_pointer == 25)
||(x_pointer == 93 && y_pointer == 25)
||(x_pointer == 94 && y_pointer == 25)
||(x_pointer == 95 && y_pointer == 25)
||(x_pointer == 96 && y_pointer == 25)
||(x_pointer == 97 && y_pointer == 25)
||(x_pointer == 98 && y_pointer == 25)
||(x_pointer == 99 && y_pointer == 25)
||(x_pointer == 100 && y_pointer == 25)
||(x_pointer == 101 && y_pointer == 25)
||(x_pointer == 102 && y_pointer == 25)
||(x_pointer == 103 && y_pointer == 25)
||(x_pointer == 104 && y_pointer == 25)
||(x_pointer == 105 && y_pointer == 25)
||(x_pointer == 106 && y_pointer == 25)
||(x_pointer == 107 && y_pointer == 25)
||(x_pointer == 108 && y_pointer == 25)
||(x_pointer == 109 && y_pointer == 25)
||(x_pointer == 110 && y_pointer == 25)
||(x_pointer == 111 && y_pointer == 25)
||(x_pointer == 112 && y_pointer == 25)
||(x_pointer == 113 && y_pointer == 25)
||(x_pointer == 114 && y_pointer == 25)
||(x_pointer == 115 && y_pointer == 25)
||(x_pointer == 116 && y_pointer == 25)
||(x_pointer == 117 && y_pointer == 25)
||(x_pointer == 43 && y_pointer == 26)
||(x_pointer == 44 && y_pointer == 26)
||(x_pointer == 45 && y_pointer == 26)
||(x_pointer == 46 && y_pointer == 26)
||(x_pointer == 47 && y_pointer == 26)
||(x_pointer == 48 && y_pointer == 26)
||(x_pointer == 49 && y_pointer == 26)
||(x_pointer == 50 && y_pointer == 26)
||(x_pointer == 51 && y_pointer == 26)
||(x_pointer == 52 && y_pointer == 26)
||(x_pointer == 53 && y_pointer == 26)
||(x_pointer == 54 && y_pointer == 26)
||(x_pointer == 55 && y_pointer == 26)
||(x_pointer == 56 && y_pointer == 26)
||(x_pointer == 57 && y_pointer == 26)
||(x_pointer == 58 && y_pointer == 26)
||(x_pointer == 59 && y_pointer == 26)
||(x_pointer == 60 && y_pointer == 26)
||(x_pointer == 61 && y_pointer == 26)
||(x_pointer == 62 && y_pointer == 26)
||(x_pointer == 63 && y_pointer == 26)
||(x_pointer == 64 && y_pointer == 26)
||(x_pointer == 65 && y_pointer == 26)
||(x_pointer == 66 && y_pointer == 26)
||(x_pointer == 67 && y_pointer == 26)
||(x_pointer == 68 && y_pointer == 26)
||(x_pointer == 69 && y_pointer == 26)
||(x_pointer == 70 && y_pointer == 26)
||(x_pointer == 90 && y_pointer == 26)
||(x_pointer == 91 && y_pointer == 26)
||(x_pointer == 92 && y_pointer == 26)
||(x_pointer == 93 && y_pointer == 26)
||(x_pointer == 94 && y_pointer == 26)
||(x_pointer == 95 && y_pointer == 26)
||(x_pointer == 96 && y_pointer == 26)
||(x_pointer == 97 && y_pointer == 26)
||(x_pointer == 98 && y_pointer == 26)
||(x_pointer == 99 && y_pointer == 26)
||(x_pointer == 100 && y_pointer == 26)
||(x_pointer == 101 && y_pointer == 26)
||(x_pointer == 102 && y_pointer == 26)
||(x_pointer == 103 && y_pointer == 26)
||(x_pointer == 104 && y_pointer == 26)
||(x_pointer == 105 && y_pointer == 26)
||(x_pointer == 106 && y_pointer == 26)
||(x_pointer == 107 && y_pointer == 26)
||(x_pointer == 108 && y_pointer == 26)
||(x_pointer == 109 && y_pointer == 26)
||(x_pointer == 110 && y_pointer == 26)
||(x_pointer == 111 && y_pointer == 26)
||(x_pointer == 112 && y_pointer == 26)
||(x_pointer == 113 && y_pointer == 26)
||(x_pointer == 114 && y_pointer == 26)
||(x_pointer == 115 && y_pointer == 26)
||(x_pointer == 116 && y_pointer == 26)
||(x_pointer == 117 && y_pointer == 26)
||(x_pointer == 43 && y_pointer == 27)
||(x_pointer == 44 && y_pointer == 27)
||(x_pointer == 45 && y_pointer == 27)
||(x_pointer == 46 && y_pointer == 27)
||(x_pointer == 47 && y_pointer == 27)
||(x_pointer == 48 && y_pointer == 27)
||(x_pointer == 49 && y_pointer == 27)
||(x_pointer == 50 && y_pointer == 27)
||(x_pointer == 51 && y_pointer == 27)
||(x_pointer == 52 && y_pointer == 27)
||(x_pointer == 53 && y_pointer == 27)
||(x_pointer == 54 && y_pointer == 27)
||(x_pointer == 55 && y_pointer == 27)
||(x_pointer == 56 && y_pointer == 27)
||(x_pointer == 57 && y_pointer == 27)
||(x_pointer == 58 && y_pointer == 27)
||(x_pointer == 59 && y_pointer == 27)
||(x_pointer == 60 && y_pointer == 27)
||(x_pointer == 61 && y_pointer == 27)
||(x_pointer == 62 && y_pointer == 27)
||(x_pointer == 63 && y_pointer == 27)
||(x_pointer == 64 && y_pointer == 27)
||(x_pointer == 65 && y_pointer == 27)
||(x_pointer == 66 && y_pointer == 27)
||(x_pointer == 67 && y_pointer == 27)
||(x_pointer == 68 && y_pointer == 27)
||(x_pointer == 69 && y_pointer == 27)
||(x_pointer == 70 && y_pointer == 27)
||(x_pointer == 90 && y_pointer == 27)
||(x_pointer == 91 && y_pointer == 27)
||(x_pointer == 92 && y_pointer == 27)
||(x_pointer == 93 && y_pointer == 27)
||(x_pointer == 94 && y_pointer == 27)
||(x_pointer == 95 && y_pointer == 27)
||(x_pointer == 96 && y_pointer == 27)
||(x_pointer == 97 && y_pointer == 27)
||(x_pointer == 98 && y_pointer == 27)
||(x_pointer == 99 && y_pointer == 27)
||(x_pointer == 100 && y_pointer == 27)
||(x_pointer == 101 && y_pointer == 27)
||(x_pointer == 102 && y_pointer == 27)
||(x_pointer == 103 && y_pointer == 27)
||(x_pointer == 104 && y_pointer == 27)
||(x_pointer == 105 && y_pointer == 27)
||(x_pointer == 106 && y_pointer == 27)
||(x_pointer == 107 && y_pointer == 27)
||(x_pointer == 108 && y_pointer == 27)
||(x_pointer == 109 && y_pointer == 27)
||(x_pointer == 110 && y_pointer == 27)
||(x_pointer == 111 && y_pointer == 27)
||(x_pointer == 112 && y_pointer == 27)
||(x_pointer == 113 && y_pointer == 27)
||(x_pointer == 114 && y_pointer == 27)
||(x_pointer == 115 && y_pointer == 27)
||(x_pointer == 116 && y_pointer == 27)
||(x_pointer == 117 && y_pointer == 27)
||(x_pointer == 43 && y_pointer == 28)
||(x_pointer == 44 && y_pointer == 28)
||(x_pointer == 45 && y_pointer == 28)
||(x_pointer == 46 && y_pointer == 28)
||(x_pointer == 47 && y_pointer == 28)
||(x_pointer == 48 && y_pointer == 28)
||(x_pointer == 49 && y_pointer == 28)
||(x_pointer == 50 && y_pointer == 28)
||(x_pointer == 51 && y_pointer == 28)
||(x_pointer == 52 && y_pointer == 28)
||(x_pointer == 53 && y_pointer == 28)
||(x_pointer == 54 && y_pointer == 28)
||(x_pointer == 55 && y_pointer == 28)
||(x_pointer == 56 && y_pointer == 28)
||(x_pointer == 57 && y_pointer == 28)
||(x_pointer == 58 && y_pointer == 28)
||(x_pointer == 59 && y_pointer == 28)
||(x_pointer == 60 && y_pointer == 28)
||(x_pointer == 61 && y_pointer == 28)
||(x_pointer == 62 && y_pointer == 28)
||(x_pointer == 63 && y_pointer == 28)
||(x_pointer == 64 && y_pointer == 28)
||(x_pointer == 65 && y_pointer == 28)
||(x_pointer == 66 && y_pointer == 28)
||(x_pointer == 67 && y_pointer == 28)
||(x_pointer == 68 && y_pointer == 28)
||(x_pointer == 69 && y_pointer == 28)
||(x_pointer == 70 && y_pointer == 28)
||(x_pointer == 90 && y_pointer == 28)
||(x_pointer == 91 && y_pointer == 28)
||(x_pointer == 92 && y_pointer == 28)
||(x_pointer == 93 && y_pointer == 28)
||(x_pointer == 94 && y_pointer == 28)
||(x_pointer == 95 && y_pointer == 28)
||(x_pointer == 96 && y_pointer == 28)
||(x_pointer == 97 && y_pointer == 28)
||(x_pointer == 98 && y_pointer == 28)
||(x_pointer == 99 && y_pointer == 28)
||(x_pointer == 100 && y_pointer == 28)
||(x_pointer == 101 && y_pointer == 28)
||(x_pointer == 102 && y_pointer == 28)
||(x_pointer == 103 && y_pointer == 28)
||(x_pointer == 104 && y_pointer == 28)
||(x_pointer == 105 && y_pointer == 28)
||(x_pointer == 106 && y_pointer == 28)
||(x_pointer == 107 && y_pointer == 28)
||(x_pointer == 108 && y_pointer == 28)
||(x_pointer == 109 && y_pointer == 28)
||(x_pointer == 110 && y_pointer == 28)
||(x_pointer == 111 && y_pointer == 28)
||(x_pointer == 112 && y_pointer == 28)
||(x_pointer == 113 && y_pointer == 28)
||(x_pointer == 114 && y_pointer == 28)
||(x_pointer == 115 && y_pointer == 28)
||(x_pointer == 116 && y_pointer == 28)
||(x_pointer == 117 && y_pointer == 28)
||(x_pointer == 43 && y_pointer == 29)
||(x_pointer == 44 && y_pointer == 29)
||(x_pointer == 45 && y_pointer == 29)
||(x_pointer == 46 && y_pointer == 29)
||(x_pointer == 47 && y_pointer == 29)
||(x_pointer == 48 && y_pointer == 29)
||(x_pointer == 49 && y_pointer == 29)
||(x_pointer == 50 && y_pointer == 29)
||(x_pointer == 51 && y_pointer == 29)
||(x_pointer == 52 && y_pointer == 29)
||(x_pointer == 53 && y_pointer == 29)
||(x_pointer == 54 && y_pointer == 29)
||(x_pointer == 55 && y_pointer == 29)
||(x_pointer == 56 && y_pointer == 29)
||(x_pointer == 57 && y_pointer == 29)
||(x_pointer == 58 && y_pointer == 29)
||(x_pointer == 59 && y_pointer == 29)
||(x_pointer == 60 && y_pointer == 29)
||(x_pointer == 61 && y_pointer == 29)
||(x_pointer == 62 && y_pointer == 29)
||(x_pointer == 63 && y_pointer == 29)
||(x_pointer == 64 && y_pointer == 29)
||(x_pointer == 65 && y_pointer == 29)
||(x_pointer == 66 && y_pointer == 29)
||(x_pointer == 67 && y_pointer == 29)
||(x_pointer == 68 && y_pointer == 29)
||(x_pointer == 69 && y_pointer == 29)
||(x_pointer == 70 && y_pointer == 29)
||(x_pointer == 90 && y_pointer == 29)
||(x_pointer == 91 && y_pointer == 29)
||(x_pointer == 92 && y_pointer == 29)
||(x_pointer == 93 && y_pointer == 29)
||(x_pointer == 94 && y_pointer == 29)
||(x_pointer == 95 && y_pointer == 29)
||(x_pointer == 96 && y_pointer == 29)
||(x_pointer == 97 && y_pointer == 29)
||(x_pointer == 98 && y_pointer == 29)
||(x_pointer == 99 && y_pointer == 29)
||(x_pointer == 100 && y_pointer == 29)
||(x_pointer == 101 && y_pointer == 29)
||(x_pointer == 102 && y_pointer == 29)
||(x_pointer == 103 && y_pointer == 29)
||(x_pointer == 104 && y_pointer == 29)
||(x_pointer == 105 && y_pointer == 29)
||(x_pointer == 106 && y_pointer == 29)
||(x_pointer == 107 && y_pointer == 29)
||(x_pointer == 108 && y_pointer == 29)
||(x_pointer == 109 && y_pointer == 29)
||(x_pointer == 110 && y_pointer == 29)
||(x_pointer == 111 && y_pointer == 29)
||(x_pointer == 112 && y_pointer == 29)
||(x_pointer == 113 && y_pointer == 29)
||(x_pointer == 114 && y_pointer == 29)
||(x_pointer == 115 && y_pointer == 29)
||(x_pointer == 116 && y_pointer == 29)
||(x_pointer == 117 && y_pointer == 29)
||(x_pointer == 43 && y_pointer == 30)
||(x_pointer == 44 && y_pointer == 30)
||(x_pointer == 45 && y_pointer == 30)
||(x_pointer == 46 && y_pointer == 30)
||(x_pointer == 47 && y_pointer == 30)
||(x_pointer == 48 && y_pointer == 30)
||(x_pointer == 49 && y_pointer == 30)
||(x_pointer == 50 && y_pointer == 30)
||(x_pointer == 51 && y_pointer == 30)
||(x_pointer == 52 && y_pointer == 30)
||(x_pointer == 53 && y_pointer == 30)
||(x_pointer == 54 && y_pointer == 30)
||(x_pointer == 55 && y_pointer == 30)
||(x_pointer == 56 && y_pointer == 30)
||(x_pointer == 57 && y_pointer == 30)
||(x_pointer == 58 && y_pointer == 30)
||(x_pointer == 59 && y_pointer == 30)
||(x_pointer == 60 && y_pointer == 30)
||(x_pointer == 61 && y_pointer == 30)
||(x_pointer == 62 && y_pointer == 30)
||(x_pointer == 63 && y_pointer == 30)
||(x_pointer == 64 && y_pointer == 30)
||(x_pointer == 65 && y_pointer == 30)
||(x_pointer == 66 && y_pointer == 30)
||(x_pointer == 67 && y_pointer == 30)
||(x_pointer == 68 && y_pointer == 30)
||(x_pointer == 69 && y_pointer == 30)
||(x_pointer == 70 && y_pointer == 30)
||(x_pointer == 90 && y_pointer == 30)
||(x_pointer == 91 && y_pointer == 30)
||(x_pointer == 92 && y_pointer == 30)
||(x_pointer == 93 && y_pointer == 30)
||(x_pointer == 94 && y_pointer == 30)
||(x_pointer == 95 && y_pointer == 30)
||(x_pointer == 96 && y_pointer == 30)
||(x_pointer == 97 && y_pointer == 30)
||(x_pointer == 98 && y_pointer == 30)
||(x_pointer == 99 && y_pointer == 30)
||(x_pointer == 100 && y_pointer == 30)
||(x_pointer == 101 && y_pointer == 30)
||(x_pointer == 102 && y_pointer == 30)
||(x_pointer == 103 && y_pointer == 30)
||(x_pointer == 104 && y_pointer == 30)
||(x_pointer == 105 && y_pointer == 30)
||(x_pointer == 106 && y_pointer == 30)
||(x_pointer == 107 && y_pointer == 30)
||(x_pointer == 108 && y_pointer == 30)
||(x_pointer == 109 && y_pointer == 30)
||(x_pointer == 110 && y_pointer == 30)
||(x_pointer == 111 && y_pointer == 30)
||(x_pointer == 112 && y_pointer == 30)
||(x_pointer == 113 && y_pointer == 30)
||(x_pointer == 114 && y_pointer == 30)
||(x_pointer == 115 && y_pointer == 30)
||(x_pointer == 116 && y_pointer == 30)
||(x_pointer == 117 && y_pointer == 30)
||(x_pointer == 43 && y_pointer == 31)
||(x_pointer == 44 && y_pointer == 31)
||(x_pointer == 45 && y_pointer == 31)
||(x_pointer == 46 && y_pointer == 31)
||(x_pointer == 47 && y_pointer == 31)
||(x_pointer == 48 && y_pointer == 31)
||(x_pointer == 49 && y_pointer == 31)
||(x_pointer == 50 && y_pointer == 31)
||(x_pointer == 51 && y_pointer == 31)
||(x_pointer == 52 && y_pointer == 31)
||(x_pointer == 53 && y_pointer == 31)
||(x_pointer == 54 && y_pointer == 31)
||(x_pointer == 55 && y_pointer == 31)
||(x_pointer == 56 && y_pointer == 31)
||(x_pointer == 57 && y_pointer == 31)
||(x_pointer == 58 && y_pointer == 31)
||(x_pointer == 59 && y_pointer == 31)
||(x_pointer == 60 && y_pointer == 31)
||(x_pointer == 61 && y_pointer == 31)
||(x_pointer == 62 && y_pointer == 31)
||(x_pointer == 63 && y_pointer == 31)
||(x_pointer == 64 && y_pointer == 31)
||(x_pointer == 65 && y_pointer == 31)
||(x_pointer == 66 && y_pointer == 31)
||(x_pointer == 67 && y_pointer == 31)
||(x_pointer == 68 && y_pointer == 31)
||(x_pointer == 69 && y_pointer == 31)
||(x_pointer == 70 && y_pointer == 31)
||(x_pointer == 90 && y_pointer == 31)
||(x_pointer == 91 && y_pointer == 31)
||(x_pointer == 92 && y_pointer == 31)
||(x_pointer == 93 && y_pointer == 31)
||(x_pointer == 94 && y_pointer == 31)
||(x_pointer == 95 && y_pointer == 31)
||(x_pointer == 96 && y_pointer == 31)
||(x_pointer == 97 && y_pointer == 31)
||(x_pointer == 98 && y_pointer == 31)
||(x_pointer == 99 && y_pointer == 31)
||(x_pointer == 100 && y_pointer == 31)
||(x_pointer == 101 && y_pointer == 31)
||(x_pointer == 102 && y_pointer == 31)
||(x_pointer == 103 && y_pointer == 31)
||(x_pointer == 104 && y_pointer == 31)
||(x_pointer == 105 && y_pointer == 31)
||(x_pointer == 106 && y_pointer == 31)
||(x_pointer == 107 && y_pointer == 31)
||(x_pointer == 108 && y_pointer == 31)
||(x_pointer == 109 && y_pointer == 31)
||(x_pointer == 110 && y_pointer == 31)
||(x_pointer == 111 && y_pointer == 31)
||(x_pointer == 112 && y_pointer == 31)
||(x_pointer == 113 && y_pointer == 31)
||(x_pointer == 114 && y_pointer == 31)
||(x_pointer == 115 && y_pointer == 31)
||(x_pointer == 116 && y_pointer == 31)
||(x_pointer == 117 && y_pointer == 31)
||(x_pointer == 43 && y_pointer == 32)
||(x_pointer == 44 && y_pointer == 32)
||(x_pointer == 45 && y_pointer == 32)
||(x_pointer == 46 && y_pointer == 32)
||(x_pointer == 47 && y_pointer == 32)
||(x_pointer == 48 && y_pointer == 32)
||(x_pointer == 49 && y_pointer == 32)
||(x_pointer == 50 && y_pointer == 32)
||(x_pointer == 51 && y_pointer == 32)
||(x_pointer == 52 && y_pointer == 32)
||(x_pointer == 53 && y_pointer == 32)
||(x_pointer == 54 && y_pointer == 32)
||(x_pointer == 55 && y_pointer == 32)
||(x_pointer == 56 && y_pointer == 32)
||(x_pointer == 57 && y_pointer == 32)
||(x_pointer == 58 && y_pointer == 32)
||(x_pointer == 59 && y_pointer == 32)
||(x_pointer == 60 && y_pointer == 32)
||(x_pointer == 61 && y_pointer == 32)
||(x_pointer == 62 && y_pointer == 32)
||(x_pointer == 63 && y_pointer == 32)
||(x_pointer == 64 && y_pointer == 32)
||(x_pointer == 65 && y_pointer == 32)
||(x_pointer == 66 && y_pointer == 32)
||(x_pointer == 67 && y_pointer == 32)
||(x_pointer == 68 && y_pointer == 32)
||(x_pointer == 69 && y_pointer == 32)
||(x_pointer == 70 && y_pointer == 32)
||(x_pointer == 90 && y_pointer == 32)
||(x_pointer == 91 && y_pointer == 32)
||(x_pointer == 92 && y_pointer == 32)
||(x_pointer == 93 && y_pointer == 32)
||(x_pointer == 94 && y_pointer == 32)
||(x_pointer == 95 && y_pointer == 32)
||(x_pointer == 96 && y_pointer == 32)
||(x_pointer == 97 && y_pointer == 32)
||(x_pointer == 98 && y_pointer == 32)
||(x_pointer == 99 && y_pointer == 32)
||(x_pointer == 100 && y_pointer == 32)
||(x_pointer == 101 && y_pointer == 32)
||(x_pointer == 102 && y_pointer == 32)
||(x_pointer == 103 && y_pointer == 32)
||(x_pointer == 104 && y_pointer == 32)
||(x_pointer == 105 && y_pointer == 32)
||(x_pointer == 106 && y_pointer == 32)
||(x_pointer == 107 && y_pointer == 32)
||(x_pointer == 108 && y_pointer == 32)
||(x_pointer == 109 && y_pointer == 32)
||(x_pointer == 110 && y_pointer == 32)
||(x_pointer == 111 && y_pointer == 32)
||(x_pointer == 112 && y_pointer == 32)
||(x_pointer == 113 && y_pointer == 32)
||(x_pointer == 114 && y_pointer == 32)
||(x_pointer == 115 && y_pointer == 32)
||(x_pointer == 116 && y_pointer == 32)
||(x_pointer == 117 && y_pointer == 32)
||(x_pointer == 43 && y_pointer == 33)
||(x_pointer == 44 && y_pointer == 33)
||(x_pointer == 45 && y_pointer == 33)
||(x_pointer == 46 && y_pointer == 33)
||(x_pointer == 47 && y_pointer == 33)
||(x_pointer == 48 && y_pointer == 33)
||(x_pointer == 49 && y_pointer == 33)
||(x_pointer == 50 && y_pointer == 33)
||(x_pointer == 51 && y_pointer == 33)
||(x_pointer == 52 && y_pointer == 33)
||(x_pointer == 53 && y_pointer == 33)
||(x_pointer == 54 && y_pointer == 33)
||(x_pointer == 55 && y_pointer == 33)
||(x_pointer == 56 && y_pointer == 33)
||(x_pointer == 57 && y_pointer == 33)
||(x_pointer == 58 && y_pointer == 33)
||(x_pointer == 59 && y_pointer == 33)
||(x_pointer == 60 && y_pointer == 33)
||(x_pointer == 61 && y_pointer == 33)
||(x_pointer == 62 && y_pointer == 33)
||(x_pointer == 63 && y_pointer == 33)
||(x_pointer == 64 && y_pointer == 33)
||(x_pointer == 65 && y_pointer == 33)
||(x_pointer == 66 && y_pointer == 33)
||(x_pointer == 67 && y_pointer == 33)
||(x_pointer == 68 && y_pointer == 33)
||(x_pointer == 69 && y_pointer == 33)
||(x_pointer == 70 && y_pointer == 33)
||(x_pointer == 90 && y_pointer == 33)
||(x_pointer == 91 && y_pointer == 33)
||(x_pointer == 92 && y_pointer == 33)
||(x_pointer == 93 && y_pointer == 33)
||(x_pointer == 94 && y_pointer == 33)
||(x_pointer == 95 && y_pointer == 33)
||(x_pointer == 96 && y_pointer == 33)
||(x_pointer == 97 && y_pointer == 33)
||(x_pointer == 98 && y_pointer == 33)
||(x_pointer == 99 && y_pointer == 33)
||(x_pointer == 100 && y_pointer == 33)
||(x_pointer == 101 && y_pointer == 33)
||(x_pointer == 102 && y_pointer == 33)
||(x_pointer == 103 && y_pointer == 33)
||(x_pointer == 104 && y_pointer == 33)
||(x_pointer == 105 && y_pointer == 33)
||(x_pointer == 106 && y_pointer == 33)
||(x_pointer == 107 && y_pointer == 33)
||(x_pointer == 108 && y_pointer == 33)
||(x_pointer == 109 && y_pointer == 33)
||(x_pointer == 110 && y_pointer == 33)
||(x_pointer == 111 && y_pointer == 33)
||(x_pointer == 112 && y_pointer == 33)
||(x_pointer == 113 && y_pointer == 33)
||(x_pointer == 114 && y_pointer == 33)
||(x_pointer == 115 && y_pointer == 33)
||(x_pointer == 116 && y_pointer == 33)
||(x_pointer == 117 && y_pointer == 33)
||(x_pointer == 43 && y_pointer == 34)
||(x_pointer == 44 && y_pointer == 34)
||(x_pointer == 45 && y_pointer == 34)
||(x_pointer == 46 && y_pointer == 34)
||(x_pointer == 47 && y_pointer == 34)
||(x_pointer == 48 && y_pointer == 34)
||(x_pointer == 49 && y_pointer == 34)
||(x_pointer == 50 && y_pointer == 34)
||(x_pointer == 51 && y_pointer == 34)
||(x_pointer == 52 && y_pointer == 34)
||(x_pointer == 53 && y_pointer == 34)
||(x_pointer == 54 && y_pointer == 34)
||(x_pointer == 55 && y_pointer == 34)
||(x_pointer == 56 && y_pointer == 34)
||(x_pointer == 57 && y_pointer == 34)
||(x_pointer == 58 && y_pointer == 34)
||(x_pointer == 59 && y_pointer == 34)
||(x_pointer == 60 && y_pointer == 34)
||(x_pointer == 61 && y_pointer == 34)
||(x_pointer == 62 && y_pointer == 34)
||(x_pointer == 63 && y_pointer == 34)
||(x_pointer == 64 && y_pointer == 34)
||(x_pointer == 65 && y_pointer == 34)
||(x_pointer == 66 && y_pointer == 34)
||(x_pointer == 67 && y_pointer == 34)
||(x_pointer == 68 && y_pointer == 34)
||(x_pointer == 69 && y_pointer == 34)
||(x_pointer == 70 && y_pointer == 34)
||(x_pointer == 90 && y_pointer == 34)
||(x_pointer == 91 && y_pointer == 34)
||(x_pointer == 92 && y_pointer == 34)
||(x_pointer == 93 && y_pointer == 34)
||(x_pointer == 94 && y_pointer == 34)
||(x_pointer == 95 && y_pointer == 34)
||(x_pointer == 96 && y_pointer == 34)
||(x_pointer == 97 && y_pointer == 34)
||(x_pointer == 98 && y_pointer == 34)
||(x_pointer == 99 && y_pointer == 34)
||(x_pointer == 100 && y_pointer == 34)
||(x_pointer == 101 && y_pointer == 34)
||(x_pointer == 102 && y_pointer == 34)
||(x_pointer == 103 && y_pointer == 34)
||(x_pointer == 104 && y_pointer == 34)
||(x_pointer == 105 && y_pointer == 34)
||(x_pointer == 106 && y_pointer == 34)
||(x_pointer == 107 && y_pointer == 34)
||(x_pointer == 108 && y_pointer == 34)
||(x_pointer == 109 && y_pointer == 34)
||(x_pointer == 110 && y_pointer == 34)
||(x_pointer == 111 && y_pointer == 34)
||(x_pointer == 112 && y_pointer == 34)
||(x_pointer == 113 && y_pointer == 34)
||(x_pointer == 114 && y_pointer == 34)
||(x_pointer == 115 && y_pointer == 34)
||(x_pointer == 116 && y_pointer == 34)
||(x_pointer == 117 && y_pointer == 34)
||(x_pointer == 43 && y_pointer == 35)
||(x_pointer == 44 && y_pointer == 35)
||(x_pointer == 45 && y_pointer == 35)
||(x_pointer == 46 && y_pointer == 35)
||(x_pointer == 47 && y_pointer == 35)
||(x_pointer == 48 && y_pointer == 35)
||(x_pointer == 49 && y_pointer == 35)
||(x_pointer == 50 && y_pointer == 35)
||(x_pointer == 51 && y_pointer == 35)
||(x_pointer == 52 && y_pointer == 35)
||(x_pointer == 53 && y_pointer == 35)
||(x_pointer == 54 && y_pointer == 35)
||(x_pointer == 55 && y_pointer == 35)
||(x_pointer == 56 && y_pointer == 35)
||(x_pointer == 57 && y_pointer == 35)
||(x_pointer == 58 && y_pointer == 35)
||(x_pointer == 59 && y_pointer == 35)
||(x_pointer == 60 && y_pointer == 35)
||(x_pointer == 61 && y_pointer == 35)
||(x_pointer == 62 && y_pointer == 35)
||(x_pointer == 63 && y_pointer == 35)
||(x_pointer == 64 && y_pointer == 35)
||(x_pointer == 65 && y_pointer == 35)
||(x_pointer == 66 && y_pointer == 35)
||(x_pointer == 67 && y_pointer == 35)
||(x_pointer == 68 && y_pointer == 35)
||(x_pointer == 69 && y_pointer == 35)
||(x_pointer == 70 && y_pointer == 35)
||(x_pointer == 90 && y_pointer == 35)
||(x_pointer == 91 && y_pointer == 35)
||(x_pointer == 92 && y_pointer == 35)
||(x_pointer == 93 && y_pointer == 35)
||(x_pointer == 94 && y_pointer == 35)
||(x_pointer == 95 && y_pointer == 35)
||(x_pointer == 96 && y_pointer == 35)
||(x_pointer == 97 && y_pointer == 35)
||(x_pointer == 98 && y_pointer == 35)
||(x_pointer == 99 && y_pointer == 35)
||(x_pointer == 100 && y_pointer == 35)
||(x_pointer == 101 && y_pointer == 35)
||(x_pointer == 102 && y_pointer == 35)
||(x_pointer == 103 && y_pointer == 35)
||(x_pointer == 104 && y_pointer == 35)
||(x_pointer == 105 && y_pointer == 35)
||(x_pointer == 106 && y_pointer == 35)
||(x_pointer == 107 && y_pointer == 35)
||(x_pointer == 108 && y_pointer == 35)
||(x_pointer == 109 && y_pointer == 35)
||(x_pointer == 110 && y_pointer == 35)
||(x_pointer == 111 && y_pointer == 35)
||(x_pointer == 112 && y_pointer == 35)
||(x_pointer == 113 && y_pointer == 35)
||(x_pointer == 114 && y_pointer == 35)
||(x_pointer == 115 && y_pointer == 35)
||(x_pointer == 116 && y_pointer == 35)
||(x_pointer == 117 && y_pointer == 35)
||(x_pointer == 43 && y_pointer == 36)
||(x_pointer == 44 && y_pointer == 36)
||(x_pointer == 45 && y_pointer == 36)
||(x_pointer == 46 && y_pointer == 36)
||(x_pointer == 47 && y_pointer == 36)
||(x_pointer == 48 && y_pointer == 36)
||(x_pointer == 49 && y_pointer == 36)
||(x_pointer == 50 && y_pointer == 36)
||(x_pointer == 51 && y_pointer == 36)
||(x_pointer == 52 && y_pointer == 36)
||(x_pointer == 53 && y_pointer == 36)
||(x_pointer == 54 && y_pointer == 36)
||(x_pointer == 55 && y_pointer == 36)
||(x_pointer == 56 && y_pointer == 36)
||(x_pointer == 57 && y_pointer == 36)
||(x_pointer == 58 && y_pointer == 36)
||(x_pointer == 59 && y_pointer == 36)
||(x_pointer == 60 && y_pointer == 36)
||(x_pointer == 61 && y_pointer == 36)
||(x_pointer == 62 && y_pointer == 36)
||(x_pointer == 63 && y_pointer == 36)
||(x_pointer == 64 && y_pointer == 36)
||(x_pointer == 65 && y_pointer == 36)
||(x_pointer == 66 && y_pointer == 36)
||(x_pointer == 67 && y_pointer == 36)
||(x_pointer == 68 && y_pointer == 36)
||(x_pointer == 69 && y_pointer == 36)
||(x_pointer == 70 && y_pointer == 36)
||(x_pointer == 90 && y_pointer == 36)
||(x_pointer == 91 && y_pointer == 36)
||(x_pointer == 92 && y_pointer == 36)
||(x_pointer == 93 && y_pointer == 36)
||(x_pointer == 94 && y_pointer == 36)
||(x_pointer == 95 && y_pointer == 36)
||(x_pointer == 96 && y_pointer == 36)
||(x_pointer == 97 && y_pointer == 36)
||(x_pointer == 98 && y_pointer == 36)
||(x_pointer == 99 && y_pointer == 36)
||(x_pointer == 100 && y_pointer == 36)
||(x_pointer == 101 && y_pointer == 36)
||(x_pointer == 102 && y_pointer == 36)
||(x_pointer == 103 && y_pointer == 36)
||(x_pointer == 104 && y_pointer == 36)
||(x_pointer == 105 && y_pointer == 36)
||(x_pointer == 106 && y_pointer == 36)
||(x_pointer == 107 && y_pointer == 36)
||(x_pointer == 108 && y_pointer == 36)
||(x_pointer == 109 && y_pointer == 36)
||(x_pointer == 110 && y_pointer == 36)
||(x_pointer == 111 && y_pointer == 36)
||(x_pointer == 112 && y_pointer == 36)
||(x_pointer == 113 && y_pointer == 36)
||(x_pointer == 114 && y_pointer == 36)
||(x_pointer == 115 && y_pointer == 36)
||(x_pointer == 116 && y_pointer == 36)
||(x_pointer == 117 && y_pointer == 36)
||(x_pointer == 43 && y_pointer == 37)
||(x_pointer == 44 && y_pointer == 37)
||(x_pointer == 45 && y_pointer == 37)
||(x_pointer == 46 && y_pointer == 37)
||(x_pointer == 47 && y_pointer == 37)
||(x_pointer == 48 && y_pointer == 37)
||(x_pointer == 49 && y_pointer == 37)
||(x_pointer == 50 && y_pointer == 37)
||(x_pointer == 51 && y_pointer == 37)
||(x_pointer == 52 && y_pointer == 37)
||(x_pointer == 53 && y_pointer == 37)
||(x_pointer == 54 && y_pointer == 37)
||(x_pointer == 55 && y_pointer == 37)
||(x_pointer == 56 && y_pointer == 37)
||(x_pointer == 57 && y_pointer == 37)
||(x_pointer == 58 && y_pointer == 37)
||(x_pointer == 59 && y_pointer == 37)
||(x_pointer == 60 && y_pointer == 37)
||(x_pointer == 61 && y_pointer == 37)
||(x_pointer == 62 && y_pointer == 37)
||(x_pointer == 63 && y_pointer == 37)
||(x_pointer == 64 && y_pointer == 37)
||(x_pointer == 65 && y_pointer == 37)
||(x_pointer == 66 && y_pointer == 37)
||(x_pointer == 67 && y_pointer == 37)
||(x_pointer == 68 && y_pointer == 37)
||(x_pointer == 69 && y_pointer == 37)
||(x_pointer == 70 && y_pointer == 37)
||(x_pointer == 90 && y_pointer == 37)
||(x_pointer == 91 && y_pointer == 37)
||(x_pointer == 92 && y_pointer == 37)
||(x_pointer == 93 && y_pointer == 37)
||(x_pointer == 94 && y_pointer == 37)
||(x_pointer == 95 && y_pointer == 37)
||(x_pointer == 96 && y_pointer == 37)
||(x_pointer == 97 && y_pointer == 37)
||(x_pointer == 98 && y_pointer == 37)
||(x_pointer == 99 && y_pointer == 37)
||(x_pointer == 100 && y_pointer == 37)
||(x_pointer == 101 && y_pointer == 37)
||(x_pointer == 102 && y_pointer == 37)
||(x_pointer == 103 && y_pointer == 37)
||(x_pointer == 104 && y_pointer == 37)
||(x_pointer == 105 && y_pointer == 37)
||(x_pointer == 106 && y_pointer == 37)
||(x_pointer == 107 && y_pointer == 37)
||(x_pointer == 108 && y_pointer == 37)
||(x_pointer == 109 && y_pointer == 37)
||(x_pointer == 110 && y_pointer == 37)
||(x_pointer == 111 && y_pointer == 37)
||(x_pointer == 112 && y_pointer == 37)
||(x_pointer == 113 && y_pointer == 37)
||(x_pointer == 114 && y_pointer == 37)
||(x_pointer == 115 && y_pointer == 37)
||(x_pointer == 116 && y_pointer == 37)
||(x_pointer == 117 && y_pointer == 37)
||(x_pointer == 43 && y_pointer == 38)
||(x_pointer == 44 && y_pointer == 38)
||(x_pointer == 45 && y_pointer == 38)
||(x_pointer == 46 && y_pointer == 38)
||(x_pointer == 47 && y_pointer == 38)
||(x_pointer == 48 && y_pointer == 38)
||(x_pointer == 49 && y_pointer == 38)
||(x_pointer == 50 && y_pointer == 38)
||(x_pointer == 51 && y_pointer == 38)
||(x_pointer == 52 && y_pointer == 38)
||(x_pointer == 53 && y_pointer == 38)
||(x_pointer == 54 && y_pointer == 38)
||(x_pointer == 55 && y_pointer == 38)
||(x_pointer == 56 && y_pointer == 38)
||(x_pointer == 57 && y_pointer == 38)
||(x_pointer == 58 && y_pointer == 38)
||(x_pointer == 59 && y_pointer == 38)
||(x_pointer == 60 && y_pointer == 38)
||(x_pointer == 61 && y_pointer == 38)
||(x_pointer == 62 && y_pointer == 38)
||(x_pointer == 63 && y_pointer == 38)
||(x_pointer == 64 && y_pointer == 38)
||(x_pointer == 65 && y_pointer == 38)
||(x_pointer == 66 && y_pointer == 38)
||(x_pointer == 67 && y_pointer == 38)
||(x_pointer == 68 && y_pointer == 38)
||(x_pointer == 69 && y_pointer == 38)
||(x_pointer == 70 && y_pointer == 38)
||(x_pointer == 90 && y_pointer == 38)
||(x_pointer == 91 && y_pointer == 38)
||(x_pointer == 92 && y_pointer == 38)
||(x_pointer == 93 && y_pointer == 38)
||(x_pointer == 94 && y_pointer == 38)
||(x_pointer == 95 && y_pointer == 38)
||(x_pointer == 96 && y_pointer == 38)
||(x_pointer == 97 && y_pointer == 38)
||(x_pointer == 98 && y_pointer == 38)
||(x_pointer == 99 && y_pointer == 38)
||(x_pointer == 100 && y_pointer == 38)
||(x_pointer == 101 && y_pointer == 38)
||(x_pointer == 102 && y_pointer == 38)
||(x_pointer == 103 && y_pointer == 38)
||(x_pointer == 104 && y_pointer == 38)
||(x_pointer == 105 && y_pointer == 38)
||(x_pointer == 106 && y_pointer == 38)
||(x_pointer == 107 && y_pointer == 38)
||(x_pointer == 108 && y_pointer == 38)
||(x_pointer == 109 && y_pointer == 38)
||(x_pointer == 110 && y_pointer == 38)
||(x_pointer == 111 && y_pointer == 38)
||(x_pointer == 112 && y_pointer == 38)
||(x_pointer == 113 && y_pointer == 38)
||(x_pointer == 114 && y_pointer == 38)
||(x_pointer == 115 && y_pointer == 38)
||(x_pointer == 116 && y_pointer == 38)
||(x_pointer == 117 && y_pointer == 38)
||(x_pointer == 43 && y_pointer == 39)
||(x_pointer == 44 && y_pointer == 39)
||(x_pointer == 45 && y_pointer == 39)
||(x_pointer == 46 && y_pointer == 39)
||(x_pointer == 47 && y_pointer == 39)
||(x_pointer == 48 && y_pointer == 39)
||(x_pointer == 49 && y_pointer == 39)
||(x_pointer == 50 && y_pointer == 39)
||(x_pointer == 51 && y_pointer == 39)
||(x_pointer == 52 && y_pointer == 39)
||(x_pointer == 53 && y_pointer == 39)
||(x_pointer == 54 && y_pointer == 39)
||(x_pointer == 55 && y_pointer == 39)
||(x_pointer == 56 && y_pointer == 39)
||(x_pointer == 57 && y_pointer == 39)
||(x_pointer == 58 && y_pointer == 39)
||(x_pointer == 59 && y_pointer == 39)
||(x_pointer == 60 && y_pointer == 39)
||(x_pointer == 61 && y_pointer == 39)
||(x_pointer == 62 && y_pointer == 39)
||(x_pointer == 63 && y_pointer == 39)
||(x_pointer == 64 && y_pointer == 39)
||(x_pointer == 65 && y_pointer == 39)
||(x_pointer == 66 && y_pointer == 39)
||(x_pointer == 67 && y_pointer == 39)
||(x_pointer == 68 && y_pointer == 39)
||(x_pointer == 69 && y_pointer == 39)
||(x_pointer == 70 && y_pointer == 39)
||(x_pointer == 90 && y_pointer == 39)
||(x_pointer == 91 && y_pointer == 39)
||(x_pointer == 92 && y_pointer == 39)
||(x_pointer == 93 && y_pointer == 39)
||(x_pointer == 94 && y_pointer == 39)
||(x_pointer == 95 && y_pointer == 39)
||(x_pointer == 96 && y_pointer == 39)
||(x_pointer == 97 && y_pointer == 39)
||(x_pointer == 98 && y_pointer == 39)
||(x_pointer == 99 && y_pointer == 39)
||(x_pointer == 100 && y_pointer == 39)
||(x_pointer == 101 && y_pointer == 39)
||(x_pointer == 102 && y_pointer == 39)
||(x_pointer == 103 && y_pointer == 39)
||(x_pointer == 104 && y_pointer == 39)
||(x_pointer == 105 && y_pointer == 39)
||(x_pointer == 106 && y_pointer == 39)
||(x_pointer == 107 && y_pointer == 39)
||(x_pointer == 108 && y_pointer == 39)
||(x_pointer == 109 && y_pointer == 39)
||(x_pointer == 110 && y_pointer == 39)
||(x_pointer == 111 && y_pointer == 39)
||(x_pointer == 112 && y_pointer == 39)
||(x_pointer == 113 && y_pointer == 39)
||(x_pointer == 114 && y_pointer == 39)
||(x_pointer == 115 && y_pointer == 39)
||(x_pointer == 116 && y_pointer == 39)
||(x_pointer == 117 && y_pointer == 39)
||(x_pointer == 43 && y_pointer == 40)
||(x_pointer == 44 && y_pointer == 40)
||(x_pointer == 45 && y_pointer == 40)
||(x_pointer == 46 && y_pointer == 40)
||(x_pointer == 47 && y_pointer == 40)
||(x_pointer == 48 && y_pointer == 40)
||(x_pointer == 49 && y_pointer == 40)
||(x_pointer == 50 && y_pointer == 40)
||(x_pointer == 51 && y_pointer == 40)
||(x_pointer == 52 && y_pointer == 40)
||(x_pointer == 53 && y_pointer == 40)
||(x_pointer == 54 && y_pointer == 40)
||(x_pointer == 55 && y_pointer == 40)
||(x_pointer == 56 && y_pointer == 40)
||(x_pointer == 57 && y_pointer == 40)
||(x_pointer == 58 && y_pointer == 40)
||(x_pointer == 59 && y_pointer == 40)
||(x_pointer == 60 && y_pointer == 40)
||(x_pointer == 61 && y_pointer == 40)
||(x_pointer == 62 && y_pointer == 40)
||(x_pointer == 63 && y_pointer == 40)
||(x_pointer == 64 && y_pointer == 40)
||(x_pointer == 65 && y_pointer == 40)
||(x_pointer == 66 && y_pointer == 40)
||(x_pointer == 67 && y_pointer == 40)
||(x_pointer == 68 && y_pointer == 40)
||(x_pointer == 69 && y_pointer == 40)
||(x_pointer == 70 && y_pointer == 40)
||(x_pointer == 90 && y_pointer == 40)
||(x_pointer == 91 && y_pointer == 40)
||(x_pointer == 92 && y_pointer == 40)
||(x_pointer == 93 && y_pointer == 40)
||(x_pointer == 94 && y_pointer == 40)
||(x_pointer == 95 && y_pointer == 40)
||(x_pointer == 96 && y_pointer == 40)
||(x_pointer == 97 && y_pointer == 40)
||(x_pointer == 98 && y_pointer == 40)
||(x_pointer == 99 && y_pointer == 40)
||(x_pointer == 100 && y_pointer == 40)
||(x_pointer == 101 && y_pointer == 40)
||(x_pointer == 102 && y_pointer == 40)
||(x_pointer == 103 && y_pointer == 40)
||(x_pointer == 104 && y_pointer == 40)
||(x_pointer == 105 && y_pointer == 40)
||(x_pointer == 106 && y_pointer == 40)
||(x_pointer == 107 && y_pointer == 40)
||(x_pointer == 108 && y_pointer == 40)
||(x_pointer == 109 && y_pointer == 40)
||(x_pointer == 110 && y_pointer == 40)
||(x_pointer == 111 && y_pointer == 40)
||(x_pointer == 112 && y_pointer == 40)
||(x_pointer == 113 && y_pointer == 40)
||(x_pointer == 114 && y_pointer == 40)
||(x_pointer == 115 && y_pointer == 40)
||(x_pointer == 116 && y_pointer == 40)
||(x_pointer == 117 && y_pointer == 40)
||(x_pointer == 43 && y_pointer == 41)
||(x_pointer == 44 && y_pointer == 41)
||(x_pointer == 45 && y_pointer == 41)
||(x_pointer == 46 && y_pointer == 41)
||(x_pointer == 47 && y_pointer == 41)
||(x_pointer == 48 && y_pointer == 41)
||(x_pointer == 49 && y_pointer == 41)
||(x_pointer == 50 && y_pointer == 41)
||(x_pointer == 51 && y_pointer == 41)
||(x_pointer == 52 && y_pointer == 41)
||(x_pointer == 53 && y_pointer == 41)
||(x_pointer == 54 && y_pointer == 41)
||(x_pointer == 55 && y_pointer == 41)
||(x_pointer == 56 && y_pointer == 41)
||(x_pointer == 57 && y_pointer == 41)
||(x_pointer == 58 && y_pointer == 41)
||(x_pointer == 59 && y_pointer == 41)
||(x_pointer == 60 && y_pointer == 41)
||(x_pointer == 61 && y_pointer == 41)
||(x_pointer == 62 && y_pointer == 41)
||(x_pointer == 63 && y_pointer == 41)
||(x_pointer == 64 && y_pointer == 41)
||(x_pointer == 65 && y_pointer == 41)
||(x_pointer == 66 && y_pointer == 41)
||(x_pointer == 67 && y_pointer == 41)
||(x_pointer == 68 && y_pointer == 41)
||(x_pointer == 69 && y_pointer == 41)
||(x_pointer == 70 && y_pointer == 41)
||(x_pointer == 90 && y_pointer == 41)
||(x_pointer == 91 && y_pointer == 41)
||(x_pointer == 92 && y_pointer == 41)
||(x_pointer == 93 && y_pointer == 41)
||(x_pointer == 94 && y_pointer == 41)
||(x_pointer == 95 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 99 && y_pointer == 41)
||(x_pointer == 100 && y_pointer == 41)
||(x_pointer == 101 && y_pointer == 41)
||(x_pointer == 102 && y_pointer == 41)
||(x_pointer == 103 && y_pointer == 41)
||(x_pointer == 104 && y_pointer == 41)
||(x_pointer == 105 && y_pointer == 41)
||(x_pointer == 106 && y_pointer == 41)
||(x_pointer == 107 && y_pointer == 41)
||(x_pointer == 108 && y_pointer == 41)
||(x_pointer == 109 && y_pointer == 41)
||(x_pointer == 110 && y_pointer == 41)
||(x_pointer == 111 && y_pointer == 41)
||(x_pointer == 112 && y_pointer == 41)
||(x_pointer == 113 && y_pointer == 41)
||(x_pointer == 114 && y_pointer == 41)
||(x_pointer == 115 && y_pointer == 41)
||(x_pointer == 116 && y_pointer == 41)
||(x_pointer == 117 && y_pointer == 41)
||(x_pointer == 43 && y_pointer == 42)
||(x_pointer == 44 && y_pointer == 42)
||(x_pointer == 45 && y_pointer == 42)
||(x_pointer == 46 && y_pointer == 42)
||(x_pointer == 47 && y_pointer == 42)
||(x_pointer == 48 && y_pointer == 42)
||(x_pointer == 49 && y_pointer == 42)
||(x_pointer == 50 && y_pointer == 42)
||(x_pointer == 51 && y_pointer == 42)
||(x_pointer == 52 && y_pointer == 42)
||(x_pointer == 53 && y_pointer == 42)
||(x_pointer == 54 && y_pointer == 42)
||(x_pointer == 55 && y_pointer == 42)
||(x_pointer == 56 && y_pointer == 42)
||(x_pointer == 57 && y_pointer == 42)
||(x_pointer == 58 && y_pointer == 42)
||(x_pointer == 59 && y_pointer == 42)
||(x_pointer == 60 && y_pointer == 42)
||(x_pointer == 61 && y_pointer == 42)
||(x_pointer == 62 && y_pointer == 42)
||(x_pointer == 63 && y_pointer == 42)
||(x_pointer == 64 && y_pointer == 42)
||(x_pointer == 65 && y_pointer == 42)
||(x_pointer == 66 && y_pointer == 42)
||(x_pointer == 67 && y_pointer == 42)
||(x_pointer == 68 && y_pointer == 42)
||(x_pointer == 69 && y_pointer == 42)
||(x_pointer == 70 && y_pointer == 42)
||(x_pointer == 90 && y_pointer == 42)
||(x_pointer == 91 && y_pointer == 42)
||(x_pointer == 92 && y_pointer == 42)
||(x_pointer == 93 && y_pointer == 42)
||(x_pointer == 94 && y_pointer == 42)
||(x_pointer == 95 && y_pointer == 42)
||(x_pointer == 96 && y_pointer == 42)
||(x_pointer == 97 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 99 && y_pointer == 42)
||(x_pointer == 100 && y_pointer == 42)
||(x_pointer == 101 && y_pointer == 42)
||(x_pointer == 102 && y_pointer == 42)
||(x_pointer == 103 && y_pointer == 42)
||(x_pointer == 104 && y_pointer == 42)
||(x_pointer == 105 && y_pointer == 42)
||(x_pointer == 106 && y_pointer == 42)
||(x_pointer == 107 && y_pointer == 42)
||(x_pointer == 108 && y_pointer == 42)
||(x_pointer == 109 && y_pointer == 42)
||(x_pointer == 110 && y_pointer == 42)
||(x_pointer == 111 && y_pointer == 42)
||(x_pointer == 112 && y_pointer == 42)
||(x_pointer == 113 && y_pointer == 42)
||(x_pointer == 114 && y_pointer == 42)
||(x_pointer == 115 && y_pointer == 42)
||(x_pointer == 116 && y_pointer == 42)
||(x_pointer == 117 && y_pointer == 42)
||(x_pointer == 43 && y_pointer == 43)
||(x_pointer == 44 && y_pointer == 43)
||(x_pointer == 45 && y_pointer == 43)
||(x_pointer == 46 && y_pointer == 43)
||(x_pointer == 47 && y_pointer == 43)
||(x_pointer == 48 && y_pointer == 43)
||(x_pointer == 49 && y_pointer == 43)
||(x_pointer == 50 && y_pointer == 43)
||(x_pointer == 51 && y_pointer == 43)
||(x_pointer == 52 && y_pointer == 43)
||(x_pointer == 53 && y_pointer == 43)
||(x_pointer == 54 && y_pointer == 43)
||(x_pointer == 55 && y_pointer == 43)
||(x_pointer == 56 && y_pointer == 43)
||(x_pointer == 57 && y_pointer == 43)
||(x_pointer == 58 && y_pointer == 43)
||(x_pointer == 59 && y_pointer == 43)
||(x_pointer == 60 && y_pointer == 43)
||(x_pointer == 61 && y_pointer == 43)
||(x_pointer == 62 && y_pointer == 43)
||(x_pointer == 63 && y_pointer == 43)
||(x_pointer == 64 && y_pointer == 43)
||(x_pointer == 65 && y_pointer == 43)
||(x_pointer == 66 && y_pointer == 43)
||(x_pointer == 67 && y_pointer == 43)
||(x_pointer == 68 && y_pointer == 43)
||(x_pointer == 69 && y_pointer == 43)
||(x_pointer == 70 && y_pointer == 43)
||(x_pointer == 90 && y_pointer == 43)
||(x_pointer == 91 && y_pointer == 43)
||(x_pointer == 92 && y_pointer == 43)
||(x_pointer == 93 && y_pointer == 43)
||(x_pointer == 94 && y_pointer == 43)
||(x_pointer == 95 && y_pointer == 43)
||(x_pointer == 96 && y_pointer == 43)
||(x_pointer == 97 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 99 && y_pointer == 43)
||(x_pointer == 100 && y_pointer == 43)
||(x_pointer == 101 && y_pointer == 43)
||(x_pointer == 102 && y_pointer == 43)
||(x_pointer == 103 && y_pointer == 43)
||(x_pointer == 104 && y_pointer == 43)
||(x_pointer == 105 && y_pointer == 43)
||(x_pointer == 106 && y_pointer == 43)
||(x_pointer == 107 && y_pointer == 43)
||(x_pointer == 108 && y_pointer == 43)
||(x_pointer == 109 && y_pointer == 43)
||(x_pointer == 110 && y_pointer == 43)
||(x_pointer == 111 && y_pointer == 43)
||(x_pointer == 112 && y_pointer == 43)
||(x_pointer == 113 && y_pointer == 43)
||(x_pointer == 114 && y_pointer == 43)
||(x_pointer == 115 && y_pointer == 43)
||(x_pointer == 116 && y_pointer == 43)
||(x_pointer == 117 && y_pointer == 43)
||(x_pointer == 43 && y_pointer == 44)
||(x_pointer == 44 && y_pointer == 44)
||(x_pointer == 45 && y_pointer == 44)
||(x_pointer == 46 && y_pointer == 44)
||(x_pointer == 47 && y_pointer == 44)
||(x_pointer == 48 && y_pointer == 44)
||(x_pointer == 49 && y_pointer == 44)
||(x_pointer == 50 && y_pointer == 44)
||(x_pointer == 51 && y_pointer == 44)
||(x_pointer == 52 && y_pointer == 44)
||(x_pointer == 53 && y_pointer == 44)
||(x_pointer == 54 && y_pointer == 44)
||(x_pointer == 55 && y_pointer == 44)
||(x_pointer == 56 && y_pointer == 44)
||(x_pointer == 57 && y_pointer == 44)
||(x_pointer == 58 && y_pointer == 44)
||(x_pointer == 59 && y_pointer == 44)
||(x_pointer == 60 && y_pointer == 44)
||(x_pointer == 61 && y_pointer == 44)
||(x_pointer == 62 && y_pointer == 44)
||(x_pointer == 63 && y_pointer == 44)
||(x_pointer == 64 && y_pointer == 44)
||(x_pointer == 65 && y_pointer == 44)
||(x_pointer == 66 && y_pointer == 44)
||(x_pointer == 67 && y_pointer == 44)
||(x_pointer == 68 && y_pointer == 44)
||(x_pointer == 69 && y_pointer == 44)
||(x_pointer == 70 && y_pointer == 44)
||(x_pointer == 90 && y_pointer == 44)
||(x_pointer == 91 && y_pointer == 44)
||(x_pointer == 92 && y_pointer == 44)
||(x_pointer == 93 && y_pointer == 44)
||(x_pointer == 94 && y_pointer == 44)
||(x_pointer == 95 && y_pointer == 44)
||(x_pointer == 96 && y_pointer == 44)
||(x_pointer == 97 && y_pointer == 44)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 99 && y_pointer == 44)
||(x_pointer == 100 && y_pointer == 44)
||(x_pointer == 101 && y_pointer == 44)
||(x_pointer == 102 && y_pointer == 44)
||(x_pointer == 103 && y_pointer == 44)
||(x_pointer == 104 && y_pointer == 44)
||(x_pointer == 105 && y_pointer == 44)
||(x_pointer == 106 && y_pointer == 44)
||(x_pointer == 107 && y_pointer == 44)
||(x_pointer == 108 && y_pointer == 44)
||(x_pointer == 109 && y_pointer == 44)
||(x_pointer == 110 && y_pointer == 44)
||(x_pointer == 111 && y_pointer == 44)
||(x_pointer == 112 && y_pointer == 44)
||(x_pointer == 113 && y_pointer == 44)
||(x_pointer == 114 && y_pointer == 44)
||(x_pointer == 115 && y_pointer == 44)
||(x_pointer == 116 && y_pointer == 44)
||(x_pointer == 117 && y_pointer == 44)
||(x_pointer == 43 && y_pointer == 45)
||(x_pointer == 44 && y_pointer == 45)
||(x_pointer == 45 && y_pointer == 45)
||(x_pointer == 46 && y_pointer == 45)
||(x_pointer == 47 && y_pointer == 45)
||(x_pointer == 48 && y_pointer == 45)
||(x_pointer == 49 && y_pointer == 45)
||(x_pointer == 50 && y_pointer == 45)
||(x_pointer == 51 && y_pointer == 45)
||(x_pointer == 52 && y_pointer == 45)
||(x_pointer == 53 && y_pointer == 45)
||(x_pointer == 54 && y_pointer == 45)
||(x_pointer == 55 && y_pointer == 45)
||(x_pointer == 56 && y_pointer == 45)
||(x_pointer == 57 && y_pointer == 45)
||(x_pointer == 58 && y_pointer == 45)
||(x_pointer == 59 && y_pointer == 45)
||(x_pointer == 60 && y_pointer == 45)
||(x_pointer == 61 && y_pointer == 45)
||(x_pointer == 62 && y_pointer == 45)
||(x_pointer == 63 && y_pointer == 45)
||(x_pointer == 64 && y_pointer == 45)
||(x_pointer == 65 && y_pointer == 45)
||(x_pointer == 66 && y_pointer == 45)
||(x_pointer == 67 && y_pointer == 45)
||(x_pointer == 68 && y_pointer == 45)
||(x_pointer == 69 && y_pointer == 45)
||(x_pointer == 70 && y_pointer == 45)
||(x_pointer == 90 && y_pointer == 45)
||(x_pointer == 91 && y_pointer == 45)
||(x_pointer == 92 && y_pointer == 45)
||(x_pointer == 93 && y_pointer == 45)
||(x_pointer == 94 && y_pointer == 45)
||(x_pointer == 95 && y_pointer == 45)
||(x_pointer == 96 && y_pointer == 45)
||(x_pointer == 97 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 99 && y_pointer == 45)
||(x_pointer == 100 && y_pointer == 45)
||(x_pointer == 101 && y_pointer == 45)
||(x_pointer == 102 && y_pointer == 45)
||(x_pointer == 103 && y_pointer == 45)
||(x_pointer == 104 && y_pointer == 45)
||(x_pointer == 105 && y_pointer == 45)
||(x_pointer == 106 && y_pointer == 45)
||(x_pointer == 107 && y_pointer == 45)
||(x_pointer == 108 && y_pointer == 45)
||(x_pointer == 109 && y_pointer == 45)
||(x_pointer == 110 && y_pointer == 45)
||(x_pointer == 111 && y_pointer == 45)
||(x_pointer == 112 && y_pointer == 45)
||(x_pointer == 113 && y_pointer == 45)
||(x_pointer == 114 && y_pointer == 45)
||(x_pointer == 115 && y_pointer == 45)
||(x_pointer == 116 && y_pointer == 45)
||(x_pointer == 117 && y_pointer == 45)
||(x_pointer == 43 && y_pointer == 46)
||(x_pointer == 44 && y_pointer == 46)
||(x_pointer == 45 && y_pointer == 46)
||(x_pointer == 46 && y_pointer == 46)
||(x_pointer == 47 && y_pointer == 46)
||(x_pointer == 48 && y_pointer == 46)
||(x_pointer == 49 && y_pointer == 46)
||(x_pointer == 50 && y_pointer == 46)
||(x_pointer == 51 && y_pointer == 46)
||(x_pointer == 52 && y_pointer == 46)
||(x_pointer == 53 && y_pointer == 46)
||(x_pointer == 54 && y_pointer == 46)
||(x_pointer == 55 && y_pointer == 46)
||(x_pointer == 56 && y_pointer == 46)
||(x_pointer == 57 && y_pointer == 46)
||(x_pointer == 58 && y_pointer == 46)
||(x_pointer == 59 && y_pointer == 46)
||(x_pointer == 60 && y_pointer == 46)
||(x_pointer == 61 && y_pointer == 46)
||(x_pointer == 62 && y_pointer == 46)
||(x_pointer == 63 && y_pointer == 46)
||(x_pointer == 64 && y_pointer == 46)
||(x_pointer == 65 && y_pointer == 46)
||(x_pointer == 66 && y_pointer == 46)
||(x_pointer == 67 && y_pointer == 46)
||(x_pointer == 68 && y_pointer == 46)
||(x_pointer == 69 && y_pointer == 46)
||(x_pointer == 70 && y_pointer == 46)
||(x_pointer == 90 && y_pointer == 46)
||(x_pointer == 91 && y_pointer == 46)
||(x_pointer == 92 && y_pointer == 46)
||(x_pointer == 93 && y_pointer == 46)
||(x_pointer == 94 && y_pointer == 46)
||(x_pointer == 95 && y_pointer == 46)
||(x_pointer == 96 && y_pointer == 46)
||(x_pointer == 97 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 99 && y_pointer == 46)
||(x_pointer == 100 && y_pointer == 46)
||(x_pointer == 101 && y_pointer == 46)
||(x_pointer == 102 && y_pointer == 46)
||(x_pointer == 103 && y_pointer == 46)
||(x_pointer == 104 && y_pointer == 46)
||(x_pointer == 105 && y_pointer == 46)
||(x_pointer == 106 && y_pointer == 46)
||(x_pointer == 107 && y_pointer == 46)
||(x_pointer == 108 && y_pointer == 46)
||(x_pointer == 109 && y_pointer == 46)
||(x_pointer == 110 && y_pointer == 46)
||(x_pointer == 111 && y_pointer == 46)
||(x_pointer == 112 && y_pointer == 46)
||(x_pointer == 113 && y_pointer == 46)
||(x_pointer == 114 && y_pointer == 46)
||(x_pointer == 115 && y_pointer == 46)
||(x_pointer == 116 && y_pointer == 46)
||(x_pointer == 117 && y_pointer == 46)
||(x_pointer == 43 && y_pointer == 47)
||(x_pointer == 44 && y_pointer == 47)
||(x_pointer == 45 && y_pointer == 47)
||(x_pointer == 46 && y_pointer == 47)
||(x_pointer == 47 && y_pointer == 47)
||(x_pointer == 48 && y_pointer == 47)
||(x_pointer == 49 && y_pointer == 47)
||(x_pointer == 50 && y_pointer == 47)
||(x_pointer == 51 && y_pointer == 47)
||(x_pointer == 52 && y_pointer == 47)
||(x_pointer == 53 && y_pointer == 47)
||(x_pointer == 54 && y_pointer == 47)
||(x_pointer == 55 && y_pointer == 47)
||(x_pointer == 56 && y_pointer == 47)
||(x_pointer == 57 && y_pointer == 47)
||(x_pointer == 58 && y_pointer == 47)
||(x_pointer == 59 && y_pointer == 47)
||(x_pointer == 60 && y_pointer == 47)
||(x_pointer == 61 && y_pointer == 47)
||(x_pointer == 62 && y_pointer == 47)
||(x_pointer == 63 && y_pointer == 47)
||(x_pointer == 64 && y_pointer == 47)
||(x_pointer == 65 && y_pointer == 47)
||(x_pointer == 66 && y_pointer == 47)
||(x_pointer == 67 && y_pointer == 47)
||(x_pointer == 68 && y_pointer == 47)
||(x_pointer == 69 && y_pointer == 47)
||(x_pointer == 70 && y_pointer == 47)
||(x_pointer == 90 && y_pointer == 47)
||(x_pointer == 91 && y_pointer == 47)
||(x_pointer == 92 && y_pointer == 47)
||(x_pointer == 93 && y_pointer == 47)
||(x_pointer == 94 && y_pointer == 47)
||(x_pointer == 95 && y_pointer == 47)
||(x_pointer == 96 && y_pointer == 47)
||(x_pointer == 97 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 99 && y_pointer == 47)
||(x_pointer == 100 && y_pointer == 47)
||(x_pointer == 101 && y_pointer == 47)
||(x_pointer == 102 && y_pointer == 47)
||(x_pointer == 103 && y_pointer == 47)
||(x_pointer == 104 && y_pointer == 47)
||(x_pointer == 105 && y_pointer == 47)
||(x_pointer == 106 && y_pointer == 47)
||(x_pointer == 107 && y_pointer == 47)
||(x_pointer == 108 && y_pointer == 47)
||(x_pointer == 109 && y_pointer == 47)
||(x_pointer == 110 && y_pointer == 47)
||(x_pointer == 111 && y_pointer == 47)
||(x_pointer == 112 && y_pointer == 47)
||(x_pointer == 113 && y_pointer == 47)
||(x_pointer == 114 && y_pointer == 47)
||(x_pointer == 115 && y_pointer == 47)
||(x_pointer == 116 && y_pointer == 47)
||(x_pointer == 117 && y_pointer == 47)
||(x_pointer == 43 && y_pointer == 48)
||(x_pointer == 44 && y_pointer == 48)
||(x_pointer == 45 && y_pointer == 48)
||(x_pointer == 46 && y_pointer == 48)
||(x_pointer == 47 && y_pointer == 48)
||(x_pointer == 48 && y_pointer == 48)
||(x_pointer == 49 && y_pointer == 48)
||(x_pointer == 50 && y_pointer == 48)
||(x_pointer == 51 && y_pointer == 48)
||(x_pointer == 52 && y_pointer == 48)
||(x_pointer == 53 && y_pointer == 48)
||(x_pointer == 54 && y_pointer == 48)
||(x_pointer == 55 && y_pointer == 48)
||(x_pointer == 56 && y_pointer == 48)
||(x_pointer == 57 && y_pointer == 48)
||(x_pointer == 58 && y_pointer == 48)
||(x_pointer == 59 && y_pointer == 48)
||(x_pointer == 60 && y_pointer == 48)
||(x_pointer == 61 && y_pointer == 48)
||(x_pointer == 62 && y_pointer == 48)
||(x_pointer == 63 && y_pointer == 48)
||(x_pointer == 64 && y_pointer == 48)
||(x_pointer == 65 && y_pointer == 48)
||(x_pointer == 66 && y_pointer == 48)
||(x_pointer == 67 && y_pointer == 48)
||(x_pointer == 68 && y_pointer == 48)
||(x_pointer == 69 && y_pointer == 48)
||(x_pointer == 70 && y_pointer == 48)
||(x_pointer == 71 && y_pointer == 48)
||(x_pointer == 72 && y_pointer == 48)
||(x_pointer == 73 && y_pointer == 48)
||(x_pointer == 74 && y_pointer == 48)
||(x_pointer == 75 && y_pointer == 48)
||(x_pointer == 76 && y_pointer == 48)
||(x_pointer == 77 && y_pointer == 48)
||(x_pointer == 78 && y_pointer == 48)
||(x_pointer == 79 && y_pointer == 48)
||(x_pointer == 80 && y_pointer == 48)
||(x_pointer == 81 && y_pointer == 48)
||(x_pointer == 82 && y_pointer == 48)
||(x_pointer == 83 && y_pointer == 48)
||(x_pointer == 84 && y_pointer == 48)
||(x_pointer == 85 && y_pointer == 48)
||(x_pointer == 86 && y_pointer == 48)
||(x_pointer == 87 && y_pointer == 48)
||(x_pointer == 88 && y_pointer == 48)
||(x_pointer == 89 && y_pointer == 48)
||(x_pointer == 90 && y_pointer == 48)
||(x_pointer == 91 && y_pointer == 48)
||(x_pointer == 92 && y_pointer == 48)
||(x_pointer == 93 && y_pointer == 48)
||(x_pointer == 94 && y_pointer == 48)
||(x_pointer == 95 && y_pointer == 48)
||(x_pointer == 96 && y_pointer == 48)
||(x_pointer == 97 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 48)
||(x_pointer == 99 && y_pointer == 48)
||(x_pointer == 100 && y_pointer == 48)
||(x_pointer == 101 && y_pointer == 48)
||(x_pointer == 102 && y_pointer == 48)
||(x_pointer == 103 && y_pointer == 48)
||(x_pointer == 104 && y_pointer == 48)
||(x_pointer == 105 && y_pointer == 48)
||(x_pointer == 106 && y_pointer == 48)
||(x_pointer == 107 && y_pointer == 48)
||(x_pointer == 108 && y_pointer == 48)
||(x_pointer == 109 && y_pointer == 48)
||(x_pointer == 110 && y_pointer == 48)
||(x_pointer == 111 && y_pointer == 48)
||(x_pointer == 112 && y_pointer == 48)
||(x_pointer == 113 && y_pointer == 48)
||(x_pointer == 114 && y_pointer == 48)
||(x_pointer == 115 && y_pointer == 48)
||(x_pointer == 116 && y_pointer == 48)
||(x_pointer == 117 && y_pointer == 48)
||(x_pointer == 70 && y_pointer == 49)
||(x_pointer == 71 && y_pointer == 49)
||(x_pointer == 72 && y_pointer == 49)
||(x_pointer == 73 && y_pointer == 49)
||(x_pointer == 74 && y_pointer == 49)
||(x_pointer == 75 && y_pointer == 49)
||(x_pointer == 76 && y_pointer == 49)
||(x_pointer == 77 && y_pointer == 49)
||(x_pointer == 78 && y_pointer == 49)
||(x_pointer == 79 && y_pointer == 49)
||(x_pointer == 80 && y_pointer == 49)
||(x_pointer == 81 && y_pointer == 49)
||(x_pointer == 82 && y_pointer == 49)
||(x_pointer == 83 && y_pointer == 49)
||(x_pointer == 84 && y_pointer == 49)
||(x_pointer == 85 && y_pointer == 49)
||(x_pointer == 86 && y_pointer == 49)
||(x_pointer == 87 && y_pointer == 49)
||(x_pointer == 88 && y_pointer == 49)
||(x_pointer == 89 && y_pointer == 49)
||(x_pointer == 90 && y_pointer == 49)
||(x_pointer == 70 && y_pointer == 50)
||(x_pointer == 71 && y_pointer == 50)
||(x_pointer == 72 && y_pointer == 50)
||(x_pointer == 73 && y_pointer == 50)
||(x_pointer == 74 && y_pointer == 50)
||(x_pointer == 75 && y_pointer == 50)
||(x_pointer == 76 && y_pointer == 50)
||(x_pointer == 77 && y_pointer == 50)
||(x_pointer == 78 && y_pointer == 50)
||(x_pointer == 79 && y_pointer == 50)
||(x_pointer == 80 && y_pointer == 50)
||(x_pointer == 81 && y_pointer == 50)
||(x_pointer == 82 && y_pointer == 50)
||(x_pointer == 83 && y_pointer == 50)
||(x_pointer == 84 && y_pointer == 50)
||(x_pointer == 85 && y_pointer == 50)
||(x_pointer == 86 && y_pointer == 50)
||(x_pointer == 87 && y_pointer == 50)
||(x_pointer == 88 && y_pointer == 50)
||(x_pointer == 89 && y_pointer == 50)
||(x_pointer == 90 && y_pointer == 50)
||(x_pointer == 70 && y_pointer == 51)
||(x_pointer == 71 && y_pointer == 51)
||(x_pointer == 72 && y_pointer == 51)
||(x_pointer == 73 && y_pointer == 51)
||(x_pointer == 74 && y_pointer == 51)
||(x_pointer == 75 && y_pointer == 51)
||(x_pointer == 76 && y_pointer == 51)
||(x_pointer == 77 && y_pointer == 51)
||(x_pointer == 78 && y_pointer == 51)
||(x_pointer == 79 && y_pointer == 51)
||(x_pointer == 80 && y_pointer == 51)
||(x_pointer == 81 && y_pointer == 51)
||(x_pointer == 82 && y_pointer == 51)
||(x_pointer == 83 && y_pointer == 51)
||(x_pointer == 84 && y_pointer == 51)
||(x_pointer == 85 && y_pointer == 51)
||(x_pointer == 86 && y_pointer == 51)
||(x_pointer == 87 && y_pointer == 51)
||(x_pointer == 88 && y_pointer == 51)
||(x_pointer == 89 && y_pointer == 51)
||(x_pointer == 90 && y_pointer == 51)
||(x_pointer == 70 && y_pointer == 52)
||(x_pointer == 71 && y_pointer == 52)
||(x_pointer == 72 && y_pointer == 52)
||(x_pointer == 73 && y_pointer == 52)
||(x_pointer == 74 && y_pointer == 52)
||(x_pointer == 75 && y_pointer == 52)
||(x_pointer == 76 && y_pointer == 52)
||(x_pointer == 77 && y_pointer == 52)
||(x_pointer == 78 && y_pointer == 52)
||(x_pointer == 79 && y_pointer == 52)
||(x_pointer == 80 && y_pointer == 52)
||(x_pointer == 81 && y_pointer == 52)
||(x_pointer == 82 && y_pointer == 52)
||(x_pointer == 83 && y_pointer == 52)
||(x_pointer == 84 && y_pointer == 52)
||(x_pointer == 85 && y_pointer == 52)
||(x_pointer == 86 && y_pointer == 52)
||(x_pointer == 87 && y_pointer == 52)
||(x_pointer == 88 && y_pointer == 52)
||(x_pointer == 89 && y_pointer == 52)
||(x_pointer == 90 && y_pointer == 52)
||(x_pointer == 70 && y_pointer == 53)
||(x_pointer == 71 && y_pointer == 53)
||(x_pointer == 72 && y_pointer == 53)
||(x_pointer == 73 && y_pointer == 53)
||(x_pointer == 74 && y_pointer == 53)
||(x_pointer == 75 && y_pointer == 53)
||(x_pointer == 76 && y_pointer == 53)
||(x_pointer == 77 && y_pointer == 53)
||(x_pointer == 78 && y_pointer == 53)
||(x_pointer == 79 && y_pointer == 53)
||(x_pointer == 80 && y_pointer == 53)
||(x_pointer == 81 && y_pointer == 53)
||(x_pointer == 82 && y_pointer == 53)
||(x_pointer == 83 && y_pointer == 53)
||(x_pointer == 84 && y_pointer == 53)
||(x_pointer == 85 && y_pointer == 53)
||(x_pointer == 86 && y_pointer == 53)
||(x_pointer == 87 && y_pointer == 53)
||(x_pointer == 88 && y_pointer == 53)
||(x_pointer == 89 && y_pointer == 53)
||(x_pointer == 90 && y_pointer == 53)
||(x_pointer == 70 && y_pointer == 54)
||(x_pointer == 71 && y_pointer == 54)
||(x_pointer == 72 && y_pointer == 54)
||(x_pointer == 73 && y_pointer == 54)
||(x_pointer == 74 && y_pointer == 54)
||(x_pointer == 75 && y_pointer == 54)
||(x_pointer == 76 && y_pointer == 54)
||(x_pointer == 77 && y_pointer == 54)
||(x_pointer == 78 && y_pointer == 54)
||(x_pointer == 79 && y_pointer == 54)
||(x_pointer == 80 && y_pointer == 54)
||(x_pointer == 81 && y_pointer == 54)
||(x_pointer == 82 && y_pointer == 54)
||(x_pointer == 83 && y_pointer == 54)
||(x_pointer == 84 && y_pointer == 54)
||(x_pointer == 85 && y_pointer == 54)
||(x_pointer == 86 && y_pointer == 54)
||(x_pointer == 87 && y_pointer == 54)
||(x_pointer == 88 && y_pointer == 54)
||(x_pointer == 89 && y_pointer == 54)
||(x_pointer == 90 && y_pointer == 54)
||(x_pointer == 70 && y_pointer == 55)
||(x_pointer == 71 && y_pointer == 55)
||(x_pointer == 72 && y_pointer == 55)
||(x_pointer == 73 && y_pointer == 55)
||(x_pointer == 74 && y_pointer == 55)
||(x_pointer == 75 && y_pointer == 55)
||(x_pointer == 76 && y_pointer == 55)
||(x_pointer == 77 && y_pointer == 55)
||(x_pointer == 78 && y_pointer == 55)
||(x_pointer == 79 && y_pointer == 55)
||(x_pointer == 80 && y_pointer == 55)
||(x_pointer == 81 && y_pointer == 55)
||(x_pointer == 82 && y_pointer == 55)
||(x_pointer == 83 && y_pointer == 55)
||(x_pointer == 84 && y_pointer == 55)
||(x_pointer == 85 && y_pointer == 55)
||(x_pointer == 86 && y_pointer == 55)
||(x_pointer == 87 && y_pointer == 55)
||(x_pointer == 88 && y_pointer == 55)
||(x_pointer == 89 && y_pointer == 55)
||(x_pointer == 90 && y_pointer == 55)
||(x_pointer == 70 && y_pointer == 56)
||(x_pointer == 71 && y_pointer == 56)
||(x_pointer == 72 && y_pointer == 56)
||(x_pointer == 73 && y_pointer == 56)
||(x_pointer == 74 && y_pointer == 56)
||(x_pointer == 75 && y_pointer == 56)
||(x_pointer == 76 && y_pointer == 56)
||(x_pointer == 77 && y_pointer == 56)
||(x_pointer == 78 && y_pointer == 56)
||(x_pointer == 79 && y_pointer == 56)
||(x_pointer == 80 && y_pointer == 56)
||(x_pointer == 81 && y_pointer == 56)
||(x_pointer == 82 && y_pointer == 56)
||(x_pointer == 83 && y_pointer == 56)
||(x_pointer == 84 && y_pointer == 56)
||(x_pointer == 85 && y_pointer == 56)
||(x_pointer == 86 && y_pointer == 56)
||(x_pointer == 87 && y_pointer == 56)
||(x_pointer == 88 && y_pointer == 56)
||(x_pointer == 89 && y_pointer == 56)
||(x_pointer == 90 && y_pointer == 56)
||(x_pointer == 70 && y_pointer == 57)
||(x_pointer == 71 && y_pointer == 57)
||(x_pointer == 72 && y_pointer == 57)
||(x_pointer == 73 && y_pointer == 57)
||(x_pointer == 74 && y_pointer == 57)
||(x_pointer == 75 && y_pointer == 57)
||(x_pointer == 76 && y_pointer == 57)
||(x_pointer == 77 && y_pointer == 57)
||(x_pointer == 78 && y_pointer == 57)
||(x_pointer == 79 && y_pointer == 57)
||(x_pointer == 80 && y_pointer == 57)
||(x_pointer == 81 && y_pointer == 57)
||(x_pointer == 82 && y_pointer == 57)
||(x_pointer == 83 && y_pointer == 57)
||(x_pointer == 84 && y_pointer == 57)
||(x_pointer == 85 && y_pointer == 57)
||(x_pointer == 86 && y_pointer == 57)
||(x_pointer == 87 && y_pointer == 57)
||(x_pointer == 88 && y_pointer == 57)
||(x_pointer == 89 && y_pointer == 57)
||(x_pointer == 90 && y_pointer == 57)
||(x_pointer == 70 && y_pointer == 58)
||(x_pointer == 71 && y_pointer == 58)
||(x_pointer == 72 && y_pointer == 58)
||(x_pointer == 73 && y_pointer == 58)
||(x_pointer == 74 && y_pointer == 58)
||(x_pointer == 75 && y_pointer == 58)
||(x_pointer == 76 && y_pointer == 58)
||(x_pointer == 77 && y_pointer == 58)
||(x_pointer == 78 && y_pointer == 58)
||(x_pointer == 79 && y_pointer == 58)
||(x_pointer == 80 && y_pointer == 58)
||(x_pointer == 81 && y_pointer == 58)
||(x_pointer == 82 && y_pointer == 58)
||(x_pointer == 83 && y_pointer == 58)
||(x_pointer == 84 && y_pointer == 58)
||(x_pointer == 85 && y_pointer == 58)
||(x_pointer == 86 && y_pointer == 58)
||(x_pointer == 87 && y_pointer == 58)
||(x_pointer == 88 && y_pointer == 58)
||(x_pointer == 89 && y_pointer == 58)
||(x_pointer == 90 && y_pointer == 58)
||(x_pointer == 70 && y_pointer == 59)
||(x_pointer == 71 && y_pointer == 59)
||(x_pointer == 72 && y_pointer == 59)
||(x_pointer == 73 && y_pointer == 59)
||(x_pointer == 74 && y_pointer == 59)
||(x_pointer == 75 && y_pointer == 59)
||(x_pointer == 76 && y_pointer == 59)
||(x_pointer == 77 && y_pointer == 59)
||(x_pointer == 78 && y_pointer == 59)
||(x_pointer == 79 && y_pointer == 59)
||(x_pointer == 80 && y_pointer == 59)
||(x_pointer == 81 && y_pointer == 59)
||(x_pointer == 82 && y_pointer == 59)
||(x_pointer == 83 && y_pointer == 59)
||(x_pointer == 84 && y_pointer == 59)
||(x_pointer == 85 && y_pointer == 59)
||(x_pointer == 86 && y_pointer == 59)
||(x_pointer == 87 && y_pointer == 59)
||(x_pointer == 88 && y_pointer == 59)
||(x_pointer == 89 && y_pointer == 59)
||(x_pointer == 90 && y_pointer == 59)
||(x_pointer == 56 && y_pointer == 60)
||(x_pointer == 57 && y_pointer == 60)
||(x_pointer == 58 && y_pointer == 60)
||(x_pointer == 59 && y_pointer == 60)
||(x_pointer == 60 && y_pointer == 60)
||(x_pointer == 61 && y_pointer == 60)
||(x_pointer == 62 && y_pointer == 60)
||(x_pointer == 63 && y_pointer == 60)
||(x_pointer == 64 && y_pointer == 60)
||(x_pointer == 65 && y_pointer == 60)
||(x_pointer == 66 && y_pointer == 60)
||(x_pointer == 67 && y_pointer == 60)
||(x_pointer == 68 && y_pointer == 60)
||(x_pointer == 69 && y_pointer == 60)
||(x_pointer == 70 && y_pointer == 60)
||(x_pointer == 71 && y_pointer == 60)
||(x_pointer == 72 && y_pointer == 60)
||(x_pointer == 73 && y_pointer == 60)
||(x_pointer == 74 && y_pointer == 60)
||(x_pointer == 75 && y_pointer == 60)
||(x_pointer == 76 && y_pointer == 60)
||(x_pointer == 77 && y_pointer == 60)
||(x_pointer == 78 && y_pointer == 60)
||(x_pointer == 79 && y_pointer == 60)
||(x_pointer == 80 && y_pointer == 60)
||(x_pointer == 81 && y_pointer == 60)
||(x_pointer == 82 && y_pointer == 60)
||(x_pointer == 83 && y_pointer == 60)
||(x_pointer == 84 && y_pointer == 60)
||(x_pointer == 85 && y_pointer == 60)
||(x_pointer == 86 && y_pointer == 60)
||(x_pointer == 87 && y_pointer == 60)
||(x_pointer == 88 && y_pointer == 60)
||(x_pointer == 89 && y_pointer == 60)
||(x_pointer == 90 && y_pointer == 60)
||(x_pointer == 91 && y_pointer == 60)
||(x_pointer == 92 && y_pointer == 60)
||(x_pointer == 93 && y_pointer == 60)
||(x_pointer == 94 && y_pointer == 60)
||(x_pointer == 95 && y_pointer == 60)
||(x_pointer == 96 && y_pointer == 60)
||(x_pointer == 97 && y_pointer == 60)
||(x_pointer == 98 && y_pointer == 60)
||(x_pointer == 99 && y_pointer == 60)
||(x_pointer == 100 && y_pointer == 60)
||(x_pointer == 101 && y_pointer == 60)
||(x_pointer == 102 && y_pointer == 60)
||(x_pointer == 103 && y_pointer == 60)
||(x_pointer == 104 && y_pointer == 60)
||(x_pointer == 56 && y_pointer == 61)
||(x_pointer == 57 && y_pointer == 61)
||(x_pointer == 58 && y_pointer == 61)
||(x_pointer == 59 && y_pointer == 61)
||(x_pointer == 60 && y_pointer == 61)
||(x_pointer == 61 && y_pointer == 61)
||(x_pointer == 62 && y_pointer == 61)
||(x_pointer == 63 && y_pointer == 61)
||(x_pointer == 64 && y_pointer == 61)
||(x_pointer == 65 && y_pointer == 61)
||(x_pointer == 66 && y_pointer == 61)
||(x_pointer == 67 && y_pointer == 61)
||(x_pointer == 68 && y_pointer == 61)
||(x_pointer == 69 && y_pointer == 61)
||(x_pointer == 70 && y_pointer == 61)
||(x_pointer == 71 && y_pointer == 61)
||(x_pointer == 72 && y_pointer == 61)
||(x_pointer == 73 && y_pointer == 61)
||(x_pointer == 74 && y_pointer == 61)
||(x_pointer == 75 && y_pointer == 61)
||(x_pointer == 76 && y_pointer == 61)
||(x_pointer == 77 && y_pointer == 61)
||(x_pointer == 78 && y_pointer == 61)
||(x_pointer == 79 && y_pointer == 61)
||(x_pointer == 80 && y_pointer == 61)
||(x_pointer == 81 && y_pointer == 61)
||(x_pointer == 82 && y_pointer == 61)
||(x_pointer == 83 && y_pointer == 61)
||(x_pointer == 84 && y_pointer == 61)
||(x_pointer == 85 && y_pointer == 61)
||(x_pointer == 86 && y_pointer == 61)
||(x_pointer == 87 && y_pointer == 61)
||(x_pointer == 88 && y_pointer == 61)
||(x_pointer == 89 && y_pointer == 61)
||(x_pointer == 90 && y_pointer == 61)
||(x_pointer == 91 && y_pointer == 61)
||(x_pointer == 92 && y_pointer == 61)
||(x_pointer == 93 && y_pointer == 61)
||(x_pointer == 94 && y_pointer == 61)
||(x_pointer == 95 && y_pointer == 61)
||(x_pointer == 96 && y_pointer == 61)
||(x_pointer == 97 && y_pointer == 61)
||(x_pointer == 98 && y_pointer == 61)
||(x_pointer == 99 && y_pointer == 61)
||(x_pointer == 100 && y_pointer == 61)
||(x_pointer == 101 && y_pointer == 61)
||(x_pointer == 102 && y_pointer == 61)
||(x_pointer == 103 && y_pointer == 61)
||(x_pointer == 104 && y_pointer == 61)
||(x_pointer == 56 && y_pointer == 62)
||(x_pointer == 57 && y_pointer == 62)
||(x_pointer == 58 && y_pointer == 62)
||(x_pointer == 59 && y_pointer == 62)
||(x_pointer == 60 && y_pointer == 62)
||(x_pointer == 61 && y_pointer == 62)
||(x_pointer == 62 && y_pointer == 62)
||(x_pointer == 63 && y_pointer == 62)
||(x_pointer == 64 && y_pointer == 62)
||(x_pointer == 65 && y_pointer == 62)
||(x_pointer == 66 && y_pointer == 62)
||(x_pointer == 67 && y_pointer == 62)
||(x_pointer == 68 && y_pointer == 62)
||(x_pointer == 69 && y_pointer == 62)
||(x_pointer == 70 && y_pointer == 62)
||(x_pointer == 71 && y_pointer == 62)
||(x_pointer == 72 && y_pointer == 62)
||(x_pointer == 73 && y_pointer == 62)
||(x_pointer == 74 && y_pointer == 62)
||(x_pointer == 75 && y_pointer == 62)
||(x_pointer == 76 && y_pointer == 62)
||(x_pointer == 77 && y_pointer == 62)
||(x_pointer == 78 && y_pointer == 62)
||(x_pointer == 79 && y_pointer == 62)
||(x_pointer == 80 && y_pointer == 62)
||(x_pointer == 81 && y_pointer == 62)
||(x_pointer == 82 && y_pointer == 62)
||(x_pointer == 83 && y_pointer == 62)
||(x_pointer == 84 && y_pointer == 62)
||(x_pointer == 85 && y_pointer == 62)
||(x_pointer == 86 && y_pointer == 62)
||(x_pointer == 87 && y_pointer == 62)
||(x_pointer == 88 && y_pointer == 62)
||(x_pointer == 89 && y_pointer == 62)
||(x_pointer == 90 && y_pointer == 62)
||(x_pointer == 91 && y_pointer == 62)
||(x_pointer == 92 && y_pointer == 62)
||(x_pointer == 93 && y_pointer == 62)
||(x_pointer == 94 && y_pointer == 62)
||(x_pointer == 95 && y_pointer == 62)
||(x_pointer == 96 && y_pointer == 62)
||(x_pointer == 97 && y_pointer == 62)
||(x_pointer == 98 && y_pointer == 62)
||(x_pointer == 99 && y_pointer == 62)
||(x_pointer == 100 && y_pointer == 62)
||(x_pointer == 101 && y_pointer == 62)
||(x_pointer == 102 && y_pointer == 62)
||(x_pointer == 103 && y_pointer == 62)
||(x_pointer == 104 && y_pointer == 62)
||(x_pointer == 56 && y_pointer == 63)
||(x_pointer == 57 && y_pointer == 63)
||(x_pointer == 58 && y_pointer == 63)
||(x_pointer == 59 && y_pointer == 63)
||(x_pointer == 60 && y_pointer == 63)
||(x_pointer == 61 && y_pointer == 63)
||(x_pointer == 62 && y_pointer == 63)
||(x_pointer == 63 && y_pointer == 63)
||(x_pointer == 64 && y_pointer == 63)
||(x_pointer == 65 && y_pointer == 63)
||(x_pointer == 66 && y_pointer == 63)
||(x_pointer == 67 && y_pointer == 63)
||(x_pointer == 68 && y_pointer == 63)
||(x_pointer == 69 && y_pointer == 63)
||(x_pointer == 70 && y_pointer == 63)
||(x_pointer == 71 && y_pointer == 63)
||(x_pointer == 72 && y_pointer == 63)
||(x_pointer == 73 && y_pointer == 63)
||(x_pointer == 74 && y_pointer == 63)
||(x_pointer == 75 && y_pointer == 63)
||(x_pointer == 76 && y_pointer == 63)
||(x_pointer == 77 && y_pointer == 63)
||(x_pointer == 78 && y_pointer == 63)
||(x_pointer == 79 && y_pointer == 63)
||(x_pointer == 80 && y_pointer == 63)
||(x_pointer == 81 && y_pointer == 63)
||(x_pointer == 82 && y_pointer == 63)
||(x_pointer == 83 && y_pointer == 63)
||(x_pointer == 84 && y_pointer == 63)
||(x_pointer == 85 && y_pointer == 63)
||(x_pointer == 86 && y_pointer == 63)
||(x_pointer == 87 && y_pointer == 63)
||(x_pointer == 88 && y_pointer == 63)
||(x_pointer == 89 && y_pointer == 63)
||(x_pointer == 90 && y_pointer == 63)
||(x_pointer == 91 && y_pointer == 63)
||(x_pointer == 92 && y_pointer == 63)
||(x_pointer == 93 && y_pointer == 63)
||(x_pointer == 94 && y_pointer == 63)
||(x_pointer == 95 && y_pointer == 63)
||(x_pointer == 96 && y_pointer == 63)
||(x_pointer == 97 && y_pointer == 63)
||(x_pointer == 98 && y_pointer == 63)
||(x_pointer == 99 && y_pointer == 63)
||(x_pointer == 100 && y_pointer == 63)
||(x_pointer == 101 && y_pointer == 63)
||(x_pointer == 102 && y_pointer == 63)
||(x_pointer == 103 && y_pointer == 63)
||(x_pointer == 104 && y_pointer == 63)
||(x_pointer == 56 && y_pointer == 64)
||(x_pointer == 57 && y_pointer == 64)
||(x_pointer == 58 && y_pointer == 64)
||(x_pointer == 59 && y_pointer == 64)
||(x_pointer == 60 && y_pointer == 64)
||(x_pointer == 61 && y_pointer == 64)
||(x_pointer == 62 && y_pointer == 64)
||(x_pointer == 63 && y_pointer == 64)
||(x_pointer == 64 && y_pointer == 64)
||(x_pointer == 65 && y_pointer == 64)
||(x_pointer == 66 && y_pointer == 64)
||(x_pointer == 67 && y_pointer == 64)
||(x_pointer == 68 && y_pointer == 64)
||(x_pointer == 69 && y_pointer == 64)
||(x_pointer == 70 && y_pointer == 64)
||(x_pointer == 71 && y_pointer == 64)
||(x_pointer == 72 && y_pointer == 64)
||(x_pointer == 73 && y_pointer == 64)
||(x_pointer == 74 && y_pointer == 64)
||(x_pointer == 75 && y_pointer == 64)
||(x_pointer == 76 && y_pointer == 64)
||(x_pointer == 77 && y_pointer == 64)
||(x_pointer == 78 && y_pointer == 64)
||(x_pointer == 79 && y_pointer == 64)
||(x_pointer == 80 && y_pointer == 64)
||(x_pointer == 81 && y_pointer == 64)
||(x_pointer == 82 && y_pointer == 64)
||(x_pointer == 83 && y_pointer == 64)
||(x_pointer == 84 && y_pointer == 64)
||(x_pointer == 85 && y_pointer == 64)
||(x_pointer == 86 && y_pointer == 64)
||(x_pointer == 87 && y_pointer == 64)
||(x_pointer == 88 && y_pointer == 64)
||(x_pointer == 89 && y_pointer == 64)
||(x_pointer == 90 && y_pointer == 64)
||(x_pointer == 91 && y_pointer == 64)
||(x_pointer == 92 && y_pointer == 64)
||(x_pointer == 93 && y_pointer == 64)
||(x_pointer == 94 && y_pointer == 64)
||(x_pointer == 95 && y_pointer == 64)
||(x_pointer == 96 && y_pointer == 64)
||(x_pointer == 97 && y_pointer == 64)
||(x_pointer == 98 && y_pointer == 64)
||(x_pointer == 99 && y_pointer == 64)
||(x_pointer == 100 && y_pointer == 64)
||(x_pointer == 101 && y_pointer == 64)
||(x_pointer == 102 && y_pointer == 64)
||(x_pointer == 103 && y_pointer == 64)
||(x_pointer == 104 && y_pointer == 64)
||(x_pointer == 56 && y_pointer == 65)
||(x_pointer == 57 && y_pointer == 65)
||(x_pointer == 58 && y_pointer == 65)
||(x_pointer == 59 && y_pointer == 65)
||(x_pointer == 60 && y_pointer == 65)
||(x_pointer == 61 && y_pointer == 65)
||(x_pointer == 62 && y_pointer == 65)
||(x_pointer == 63 && y_pointer == 65)
||(x_pointer == 64 && y_pointer == 65)
||(x_pointer == 65 && y_pointer == 65)
||(x_pointer == 66 && y_pointer == 65)
||(x_pointer == 67 && y_pointer == 65)
||(x_pointer == 68 && y_pointer == 65)
||(x_pointer == 69 && y_pointer == 65)
||(x_pointer == 70 && y_pointer == 65)
||(x_pointer == 71 && y_pointer == 65)
||(x_pointer == 72 && y_pointer == 65)
||(x_pointer == 73 && y_pointer == 65)
||(x_pointer == 74 && y_pointer == 65)
||(x_pointer == 75 && y_pointer == 65)
||(x_pointer == 76 && y_pointer == 65)
||(x_pointer == 77 && y_pointer == 65)
||(x_pointer == 78 && y_pointer == 65)
||(x_pointer == 79 && y_pointer == 65)
||(x_pointer == 80 && y_pointer == 65)
||(x_pointer == 81 && y_pointer == 65)
||(x_pointer == 82 && y_pointer == 65)
||(x_pointer == 83 && y_pointer == 65)
||(x_pointer == 84 && y_pointer == 65)
||(x_pointer == 85 && y_pointer == 65)
||(x_pointer == 86 && y_pointer == 65)
||(x_pointer == 87 && y_pointer == 65)
||(x_pointer == 88 && y_pointer == 65)
||(x_pointer == 89 && y_pointer == 65)
||(x_pointer == 90 && y_pointer == 65)
||(x_pointer == 91 && y_pointer == 65)
||(x_pointer == 92 && y_pointer == 65)
||(x_pointer == 93 && y_pointer == 65)
||(x_pointer == 94 && y_pointer == 65)
||(x_pointer == 95 && y_pointer == 65)
||(x_pointer == 96 && y_pointer == 65)
||(x_pointer == 97 && y_pointer == 65)
||(x_pointer == 98 && y_pointer == 65)
||(x_pointer == 99 && y_pointer == 65)
||(x_pointer == 100 && y_pointer == 65)
||(x_pointer == 101 && y_pointer == 65)
||(x_pointer == 102 && y_pointer == 65)
||(x_pointer == 103 && y_pointer == 65)
||(x_pointer == 104 && y_pointer == 65)
||(x_pointer == 56 && y_pointer == 66)
||(x_pointer == 57 && y_pointer == 66)
||(x_pointer == 58 && y_pointer == 66)
||(x_pointer == 59 && y_pointer == 66)
||(x_pointer == 60 && y_pointer == 66)
||(x_pointer == 61 && y_pointer == 66)
||(x_pointer == 62 && y_pointer == 66)
||(x_pointer == 63 && y_pointer == 66)
||(x_pointer == 64 && y_pointer == 66)
||(x_pointer == 65 && y_pointer == 66)
||(x_pointer == 66 && y_pointer == 66)
||(x_pointer == 67 && y_pointer == 66)
||(x_pointer == 68 && y_pointer == 66)
||(x_pointer == 69 && y_pointer == 66)
||(x_pointer == 70 && y_pointer == 66)
||(x_pointer == 71 && y_pointer == 66)
||(x_pointer == 72 && y_pointer == 66)
||(x_pointer == 73 && y_pointer == 66)
||(x_pointer == 74 && y_pointer == 66)
||(x_pointer == 75 && y_pointer == 66)
||(x_pointer == 76 && y_pointer == 66)
||(x_pointer == 77 && y_pointer == 66)
||(x_pointer == 78 && y_pointer == 66)
||(x_pointer == 79 && y_pointer == 66)
||(x_pointer == 80 && y_pointer == 66)
||(x_pointer == 81 && y_pointer == 66)
||(x_pointer == 82 && y_pointer == 66)
||(x_pointer == 83 && y_pointer == 66)
||(x_pointer == 84 && y_pointer == 66)
||(x_pointer == 85 && y_pointer == 66)
||(x_pointer == 86 && y_pointer == 66)
||(x_pointer == 87 && y_pointer == 66)
||(x_pointer == 88 && y_pointer == 66)
||(x_pointer == 89 && y_pointer == 66)
||(x_pointer == 90 && y_pointer == 66)
||(x_pointer == 91 && y_pointer == 66)
||(x_pointer == 92 && y_pointer == 66)
||(x_pointer == 93 && y_pointer == 66)
||(x_pointer == 94 && y_pointer == 66)
||(x_pointer == 95 && y_pointer == 66)
||(x_pointer == 96 && y_pointer == 66)
||(x_pointer == 97 && y_pointer == 66)
||(x_pointer == 98 && y_pointer == 66)
||(x_pointer == 99 && y_pointer == 66)
||(x_pointer == 100 && y_pointer == 66)
||(x_pointer == 101 && y_pointer == 66)
||(x_pointer == 102 && y_pointer == 66)
||(x_pointer == 103 && y_pointer == 66)
||(x_pointer == 104 && y_pointer == 66)
||(x_pointer == 56 && y_pointer == 67)
||(x_pointer == 57 && y_pointer == 67)
||(x_pointer == 58 && y_pointer == 67)
||(x_pointer == 59 && y_pointer == 67)
||(x_pointer == 60 && y_pointer == 67)
||(x_pointer == 61 && y_pointer == 67)
||(x_pointer == 62 && y_pointer == 67)
||(x_pointer == 63 && y_pointer == 67)
||(x_pointer == 64 && y_pointer == 67)
||(x_pointer == 65 && y_pointer == 67)
||(x_pointer == 66 && y_pointer == 67)
||(x_pointer == 67 && y_pointer == 67)
||(x_pointer == 68 && y_pointer == 67)
||(x_pointer == 69 && y_pointer == 67)
||(x_pointer == 70 && y_pointer == 67)
||(x_pointer == 71 && y_pointer == 67)
||(x_pointer == 72 && y_pointer == 67)
||(x_pointer == 73 && y_pointer == 67)
||(x_pointer == 74 && y_pointer == 67)
||(x_pointer == 75 && y_pointer == 67)
||(x_pointer == 76 && y_pointer == 67)
||(x_pointer == 77 && y_pointer == 67)
||(x_pointer == 78 && y_pointer == 67)
||(x_pointer == 79 && y_pointer == 67)
||(x_pointer == 80 && y_pointer == 67)
||(x_pointer == 81 && y_pointer == 67)
||(x_pointer == 82 && y_pointer == 67)
||(x_pointer == 83 && y_pointer == 67)
||(x_pointer == 84 && y_pointer == 67)
||(x_pointer == 85 && y_pointer == 67)
||(x_pointer == 86 && y_pointer == 67)
||(x_pointer == 87 && y_pointer == 67)
||(x_pointer == 88 && y_pointer == 67)
||(x_pointer == 89 && y_pointer == 67)
||(x_pointer == 90 && y_pointer == 67)
||(x_pointer == 91 && y_pointer == 67)
||(x_pointer == 92 && y_pointer == 67)
||(x_pointer == 93 && y_pointer == 67)
||(x_pointer == 94 && y_pointer == 67)
||(x_pointer == 95 && y_pointer == 67)
||(x_pointer == 96 && y_pointer == 67)
||(x_pointer == 97 && y_pointer == 67)
||(x_pointer == 98 && y_pointer == 67)
||(x_pointer == 99 && y_pointer == 67)
||(x_pointer == 100 && y_pointer == 67)
||(x_pointer == 101 && y_pointer == 67)
||(x_pointer == 102 && y_pointer == 67)
||(x_pointer == 103 && y_pointer == 67)
||(x_pointer == 104 && y_pointer == 67)
||(x_pointer == 56 && y_pointer == 68)
||(x_pointer == 57 && y_pointer == 68)
||(x_pointer == 58 && y_pointer == 68)
||(x_pointer == 59 && y_pointer == 68)
||(x_pointer == 60 && y_pointer == 68)
||(x_pointer == 61 && y_pointer == 68)
||(x_pointer == 62 && y_pointer == 68)
||(x_pointer == 63 && y_pointer == 68)
||(x_pointer == 64 && y_pointer == 68)
||(x_pointer == 65 && y_pointer == 68)
||(x_pointer == 66 && y_pointer == 68)
||(x_pointer == 67 && y_pointer == 68)
||(x_pointer == 68 && y_pointer == 68)
||(x_pointer == 69 && y_pointer == 68)
||(x_pointer == 70 && y_pointer == 68)
||(x_pointer == 71 && y_pointer == 68)
||(x_pointer == 72 && y_pointer == 68)
||(x_pointer == 73 && y_pointer == 68)
||(x_pointer == 74 && y_pointer == 68)
||(x_pointer == 75 && y_pointer == 68)
||(x_pointer == 76 && y_pointer == 68)
||(x_pointer == 77 && y_pointer == 68)
||(x_pointer == 78 && y_pointer == 68)
||(x_pointer == 79 && y_pointer == 68)
||(x_pointer == 80 && y_pointer == 68)
||(x_pointer == 81 && y_pointer == 68)
||(x_pointer == 82 && y_pointer == 68)
||(x_pointer == 83 && y_pointer == 68)
||(x_pointer == 84 && y_pointer == 68)
||(x_pointer == 85 && y_pointer == 68)
||(x_pointer == 86 && y_pointer == 68)
||(x_pointer == 87 && y_pointer == 68)
||(x_pointer == 88 && y_pointer == 68)
||(x_pointer == 89 && y_pointer == 68)
||(x_pointer == 90 && y_pointer == 68)
||(x_pointer == 91 && y_pointer == 68)
||(x_pointer == 92 && y_pointer == 68)
||(x_pointer == 93 && y_pointer == 68)
||(x_pointer == 94 && y_pointer == 68)
||(x_pointer == 95 && y_pointer == 68)
||(x_pointer == 96 && y_pointer == 68)
||(x_pointer == 97 && y_pointer == 68)
||(x_pointer == 98 && y_pointer == 68)
||(x_pointer == 99 && y_pointer == 68)
||(x_pointer == 100 && y_pointer == 68)
||(x_pointer == 101 && y_pointer == 68)
||(x_pointer == 102 && y_pointer == 68)
||(x_pointer == 103 && y_pointer == 68)
||(x_pointer == 104 && y_pointer == 68)
||(x_pointer == 56 && y_pointer == 69)
||(x_pointer == 57 && y_pointer == 69)
||(x_pointer == 58 && y_pointer == 69)
||(x_pointer == 59 && y_pointer == 69)
||(x_pointer == 60 && y_pointer == 69)
||(x_pointer == 61 && y_pointer == 69)
||(x_pointer == 62 && y_pointer == 69)
||(x_pointer == 63 && y_pointer == 69)
||(x_pointer == 64 && y_pointer == 69)
||(x_pointer == 65 && y_pointer == 69)
||(x_pointer == 66 && y_pointer == 69)
||(x_pointer == 67 && y_pointer == 69)
||(x_pointer == 68 && y_pointer == 69)
||(x_pointer == 69 && y_pointer == 69)
||(x_pointer == 70 && y_pointer == 69)
||(x_pointer == 71 && y_pointer == 69)
||(x_pointer == 72 && y_pointer == 69)
||(x_pointer == 73 && y_pointer == 69)
||(x_pointer == 74 && y_pointer == 69)
||(x_pointer == 75 && y_pointer == 69)
||(x_pointer == 76 && y_pointer == 69)
||(x_pointer == 77 && y_pointer == 69)
||(x_pointer == 78 && y_pointer == 69)
||(x_pointer == 79 && y_pointer == 69)
||(x_pointer == 80 && y_pointer == 69)
||(x_pointer == 81 && y_pointer == 69)
||(x_pointer == 82 && y_pointer == 69)
||(x_pointer == 83 && y_pointer == 69)
||(x_pointer == 84 && y_pointer == 69)
||(x_pointer == 85 && y_pointer == 69)
||(x_pointer == 86 && y_pointer == 69)
||(x_pointer == 87 && y_pointer == 69)
||(x_pointer == 88 && y_pointer == 69)
||(x_pointer == 89 && y_pointer == 69)
||(x_pointer == 90 && y_pointer == 69)
||(x_pointer == 91 && y_pointer == 69)
||(x_pointer == 92 && y_pointer == 69)
||(x_pointer == 93 && y_pointer == 69)
||(x_pointer == 94 && y_pointer == 69)
||(x_pointer == 95 && y_pointer == 69)
||(x_pointer == 96 && y_pointer == 69)
||(x_pointer == 97 && y_pointer == 69)
||(x_pointer == 98 && y_pointer == 69)
||(x_pointer == 99 && y_pointer == 69)
||(x_pointer == 100 && y_pointer == 69)
||(x_pointer == 101 && y_pointer == 69)
||(x_pointer == 102 && y_pointer == 69)
||(x_pointer == 103 && y_pointer == 69)
||(x_pointer == 104 && y_pointer == 69)
||(x_pointer == 56 && y_pointer == 70)
||(x_pointer == 57 && y_pointer == 70)
||(x_pointer == 58 && y_pointer == 70)
||(x_pointer == 59 && y_pointer == 70)
||(x_pointer == 60 && y_pointer == 70)
||(x_pointer == 61 && y_pointer == 70)
||(x_pointer == 62 && y_pointer == 70)
||(x_pointer == 63 && y_pointer == 70)
||(x_pointer == 64 && y_pointer == 70)
||(x_pointer == 65 && y_pointer == 70)
||(x_pointer == 66 && y_pointer == 70)
||(x_pointer == 67 && y_pointer == 70)
||(x_pointer == 68 && y_pointer == 70)
||(x_pointer == 69 && y_pointer == 70)
||(x_pointer == 70 && y_pointer == 70)
||(x_pointer == 71 && y_pointer == 70)
||(x_pointer == 72 && y_pointer == 70)
||(x_pointer == 73 && y_pointer == 70)
||(x_pointer == 74 && y_pointer == 70)
||(x_pointer == 75 && y_pointer == 70)
||(x_pointer == 76 && y_pointer == 70)
||(x_pointer == 77 && y_pointer == 70)
||(x_pointer == 78 && y_pointer == 70)
||(x_pointer == 79 && y_pointer == 70)
||(x_pointer == 80 && y_pointer == 70)
||(x_pointer == 81 && y_pointer == 70)
||(x_pointer == 82 && y_pointer == 70)
||(x_pointer == 83 && y_pointer == 70)
||(x_pointer == 84 && y_pointer == 70)
||(x_pointer == 85 && y_pointer == 70)
||(x_pointer == 86 && y_pointer == 70)
||(x_pointer == 87 && y_pointer == 70)
||(x_pointer == 88 && y_pointer == 70)
||(x_pointer == 89 && y_pointer == 70)
||(x_pointer == 90 && y_pointer == 70)
||(x_pointer == 91 && y_pointer == 70)
||(x_pointer == 92 && y_pointer == 70)
||(x_pointer == 93 && y_pointer == 70)
||(x_pointer == 94 && y_pointer == 70)
||(x_pointer == 95 && y_pointer == 70)
||(x_pointer == 96 && y_pointer == 70)
||(x_pointer == 97 && y_pointer == 70)
||(x_pointer == 98 && y_pointer == 70)
||(x_pointer == 99 && y_pointer == 70)
||(x_pointer == 100 && y_pointer == 70)
||(x_pointer == 101 && y_pointer == 70)
||(x_pointer == 102 && y_pointer == 70)
||(x_pointer == 103 && y_pointer == 70)
||(x_pointer == 104 && y_pointer == 70)
||(x_pointer == 56 && y_pointer == 71)
||(x_pointer == 57 && y_pointer == 71)
||(x_pointer == 58 && y_pointer == 71)
||(x_pointer == 59 && y_pointer == 71)
||(x_pointer == 60 && y_pointer == 71)
||(x_pointer == 61 && y_pointer == 71)
||(x_pointer == 62 && y_pointer == 71)
||(x_pointer == 63 && y_pointer == 71)
||(x_pointer == 64 && y_pointer == 71)
||(x_pointer == 65 && y_pointer == 71)
||(x_pointer == 66 && y_pointer == 71)
||(x_pointer == 67 && y_pointer == 71)
||(x_pointer == 68 && y_pointer == 71)
||(x_pointer == 69 && y_pointer == 71)
||(x_pointer == 70 && y_pointer == 71)
||(x_pointer == 71 && y_pointer == 71)
||(x_pointer == 72 && y_pointer == 71)
||(x_pointer == 73 && y_pointer == 71)
||(x_pointer == 74 && y_pointer == 71)
||(x_pointer == 75 && y_pointer == 71)
||(x_pointer == 76 && y_pointer == 71)
||(x_pointer == 77 && y_pointer == 71)
||(x_pointer == 78 && y_pointer == 71)
||(x_pointer == 79 && y_pointer == 71)
||(x_pointer == 80 && y_pointer == 71)
||(x_pointer == 81 && y_pointer == 71)
||(x_pointer == 82 && y_pointer == 71)
||(x_pointer == 83 && y_pointer == 71)
||(x_pointer == 84 && y_pointer == 71)
||(x_pointer == 85 && y_pointer == 71)
||(x_pointer == 86 && y_pointer == 71)
||(x_pointer == 87 && y_pointer == 71)
||(x_pointer == 88 && y_pointer == 71)
||(x_pointer == 89 && y_pointer == 71)
||(x_pointer == 90 && y_pointer == 71)
||(x_pointer == 91 && y_pointer == 71)
||(x_pointer == 92 && y_pointer == 71)
||(x_pointer == 93 && y_pointer == 71)
||(x_pointer == 94 && y_pointer == 71)
||(x_pointer == 95 && y_pointer == 71)
||(x_pointer == 96 && y_pointer == 71)
||(x_pointer == 97 && y_pointer == 71)
||(x_pointer == 98 && y_pointer == 71)
||(x_pointer == 99 && y_pointer == 71)
||(x_pointer == 100 && y_pointer == 71)
||(x_pointer == 101 && y_pointer == 71)
||(x_pointer == 102 && y_pointer == 71)
||(x_pointer == 103 && y_pointer == 71)
||(x_pointer == 104 && y_pointer == 71)
||(x_pointer == 56 && y_pointer == 72)
||(x_pointer == 57 && y_pointer == 72)
||(x_pointer == 58 && y_pointer == 72)
||(x_pointer == 59 && y_pointer == 72)
||(x_pointer == 60 && y_pointer == 72)
||(x_pointer == 61 && y_pointer == 72)
||(x_pointer == 62 && y_pointer == 72)
||(x_pointer == 63 && y_pointer == 72)
||(x_pointer == 64 && y_pointer == 72)
||(x_pointer == 65 && y_pointer == 72)
||(x_pointer == 66 && y_pointer == 72)
||(x_pointer == 67 && y_pointer == 72)
||(x_pointer == 68 && y_pointer == 72)
||(x_pointer == 69 && y_pointer == 72)
||(x_pointer == 70 && y_pointer == 72)
||(x_pointer == 71 && y_pointer == 72)
||(x_pointer == 72 && y_pointer == 72)
||(x_pointer == 73 && y_pointer == 72)
||(x_pointer == 74 && y_pointer == 72)
||(x_pointer == 75 && y_pointer == 72)
||(x_pointer == 76 && y_pointer == 72)
||(x_pointer == 77 && y_pointer == 72)
||(x_pointer == 78 && y_pointer == 72)
||(x_pointer == 79 && y_pointer == 72)
||(x_pointer == 80 && y_pointer == 72)
||(x_pointer == 81 && y_pointer == 72)
||(x_pointer == 82 && y_pointer == 72)
||(x_pointer == 83 && y_pointer == 72)
||(x_pointer == 84 && y_pointer == 72)
||(x_pointer == 85 && y_pointer == 72)
||(x_pointer == 86 && y_pointer == 72)
||(x_pointer == 87 && y_pointer == 72)
||(x_pointer == 88 && y_pointer == 72)
||(x_pointer == 89 && y_pointer == 72)
||(x_pointer == 90 && y_pointer == 72)
||(x_pointer == 91 && y_pointer == 72)
||(x_pointer == 92 && y_pointer == 72)
||(x_pointer == 93 && y_pointer == 72)
||(x_pointer == 94 && y_pointer == 72)
||(x_pointer == 95 && y_pointer == 72)
||(x_pointer == 96 && y_pointer == 72)
||(x_pointer == 97 && y_pointer == 72)
||(x_pointer == 98 && y_pointer == 72)
||(x_pointer == 99 && y_pointer == 72)
||(x_pointer == 100 && y_pointer == 72)
||(x_pointer == 101 && y_pointer == 72)
||(x_pointer == 102 && y_pointer == 72)
||(x_pointer == 103 && y_pointer == 72)
||(x_pointer == 104 && y_pointer == 72)
||(x_pointer == 56 && y_pointer == 73)
||(x_pointer == 57 && y_pointer == 73)
||(x_pointer == 58 && y_pointer == 73)
||(x_pointer == 59 && y_pointer == 73)
||(x_pointer == 60 && y_pointer == 73)
||(x_pointer == 61 && y_pointer == 73)
||(x_pointer == 62 && y_pointer == 73)
||(x_pointer == 63 && y_pointer == 73)
||(x_pointer == 64 && y_pointer == 73)
||(x_pointer == 65 && y_pointer == 73)
||(x_pointer == 66 && y_pointer == 73)
||(x_pointer == 67 && y_pointer == 73)
||(x_pointer == 68 && y_pointer == 73)
||(x_pointer == 69 && y_pointer == 73)
||(x_pointer == 70 && y_pointer == 73)
||(x_pointer == 71 && y_pointer == 73)
||(x_pointer == 72 && y_pointer == 73)
||(x_pointer == 73 && y_pointer == 73)
||(x_pointer == 74 && y_pointer == 73)
||(x_pointer == 75 && y_pointer == 73)
||(x_pointer == 76 && y_pointer == 73)
||(x_pointer == 77 && y_pointer == 73)
||(x_pointer == 78 && y_pointer == 73)
||(x_pointer == 79 && y_pointer == 73)
||(x_pointer == 80 && y_pointer == 73)
||(x_pointer == 81 && y_pointer == 73)
||(x_pointer == 82 && y_pointer == 73)
||(x_pointer == 83 && y_pointer == 73)
||(x_pointer == 84 && y_pointer == 73)
||(x_pointer == 85 && y_pointer == 73)
||(x_pointer == 86 && y_pointer == 73)
||(x_pointer == 87 && y_pointer == 73)
||(x_pointer == 88 && y_pointer == 73)
||(x_pointer == 89 && y_pointer == 73)
||(x_pointer == 90 && y_pointer == 73)
||(x_pointer == 91 && y_pointer == 73)
||(x_pointer == 92 && y_pointer == 73)
||(x_pointer == 93 && y_pointer == 73)
||(x_pointer == 94 && y_pointer == 73)
||(x_pointer == 95 && y_pointer == 73)
||(x_pointer == 96 && y_pointer == 73)
||(x_pointer == 97 && y_pointer == 73)
||(x_pointer == 98 && y_pointer == 73)
||(x_pointer == 99 && y_pointer == 73)
||(x_pointer == 100 && y_pointer == 73)
||(x_pointer == 101 && y_pointer == 73)
||(x_pointer == 102 && y_pointer == 73)
||(x_pointer == 103 && y_pointer == 73)
||(x_pointer == 104 && y_pointer == 73)
||(x_pointer == 56 && y_pointer == 74)
||(x_pointer == 57 && y_pointer == 74)
||(x_pointer == 58 && y_pointer == 74)
||(x_pointer == 59 && y_pointer == 74)
||(x_pointer == 60 && y_pointer == 74)
||(x_pointer == 61 && y_pointer == 74)
||(x_pointer == 62 && y_pointer == 74)
||(x_pointer == 63 && y_pointer == 74)
||(x_pointer == 64 && y_pointer == 74)
||(x_pointer == 65 && y_pointer == 74)
||(x_pointer == 66 && y_pointer == 74)
||(x_pointer == 67 && y_pointer == 74)
||(x_pointer == 68 && y_pointer == 74)
||(x_pointer == 69 && y_pointer == 74)
||(x_pointer == 70 && y_pointer == 74)
||(x_pointer == 71 && y_pointer == 74)
||(x_pointer == 72 && y_pointer == 74)
||(x_pointer == 73 && y_pointer == 74)
||(x_pointer == 74 && y_pointer == 74)
||(x_pointer == 75 && y_pointer == 74)
||(x_pointer == 76 && y_pointer == 74)
||(x_pointer == 77 && y_pointer == 74)
||(x_pointer == 78 && y_pointer == 74)
||(x_pointer == 79 && y_pointer == 74)
||(x_pointer == 80 && y_pointer == 74)
||(x_pointer == 81 && y_pointer == 74)
||(x_pointer == 82 && y_pointer == 74)
||(x_pointer == 83 && y_pointer == 74)
||(x_pointer == 84 && y_pointer == 74)
||(x_pointer == 85 && y_pointer == 74)
||(x_pointer == 86 && y_pointer == 74)
||(x_pointer == 87 && y_pointer == 74)
||(x_pointer == 88 && y_pointer == 74)
||(x_pointer == 89 && y_pointer == 74)
||(x_pointer == 90 && y_pointer == 74)
||(x_pointer == 91 && y_pointer == 74)
||(x_pointer == 92 && y_pointer == 74)
||(x_pointer == 93 && y_pointer == 74)
||(x_pointer == 94 && y_pointer == 74)
||(x_pointer == 95 && y_pointer == 74)
||(x_pointer == 96 && y_pointer == 74)
||(x_pointer == 97 && y_pointer == 74)
||(x_pointer == 98 && y_pointer == 74)
||(x_pointer == 99 && y_pointer == 74)
||(x_pointer == 100 && y_pointer == 74)
||(x_pointer == 101 && y_pointer == 74)
||(x_pointer == 102 && y_pointer == 74)
||(x_pointer == 103 && y_pointer == 74)
||(x_pointer == 104 && y_pointer == 74)
||(x_pointer == 56 && y_pointer == 75)
||(x_pointer == 57 && y_pointer == 75)
||(x_pointer == 58 && y_pointer == 75)
||(x_pointer == 59 && y_pointer == 75)
||(x_pointer == 60 && y_pointer == 75)
||(x_pointer == 61 && y_pointer == 75)
||(x_pointer == 62 && y_pointer == 75)
||(x_pointer == 63 && y_pointer == 75)
||(x_pointer == 64 && y_pointer == 75)
||(x_pointer == 65 && y_pointer == 75)
||(x_pointer == 66 && y_pointer == 75)
||(x_pointer == 67 && y_pointer == 75)
||(x_pointer == 68 && y_pointer == 75)
||(x_pointer == 69 && y_pointer == 75)
||(x_pointer == 70 && y_pointer == 75)
||(x_pointer == 71 && y_pointer == 75)
||(x_pointer == 72 && y_pointer == 75)
||(x_pointer == 73 && y_pointer == 75)
||(x_pointer == 74 && y_pointer == 75)
||(x_pointer == 75 && y_pointer == 75)
||(x_pointer == 76 && y_pointer == 75)
||(x_pointer == 77 && y_pointer == 75)
||(x_pointer == 78 && y_pointer == 75)
||(x_pointer == 79 && y_pointer == 75)
||(x_pointer == 80 && y_pointer == 75)
||(x_pointer == 81 && y_pointer == 75)
||(x_pointer == 82 && y_pointer == 75)
||(x_pointer == 83 && y_pointer == 75)
||(x_pointer == 84 && y_pointer == 75)
||(x_pointer == 85 && y_pointer == 75)
||(x_pointer == 86 && y_pointer == 75)
||(x_pointer == 87 && y_pointer == 75)
||(x_pointer == 88 && y_pointer == 75)
||(x_pointer == 89 && y_pointer == 75)
||(x_pointer == 90 && y_pointer == 75)
||(x_pointer == 91 && y_pointer == 75)
||(x_pointer == 92 && y_pointer == 75)
||(x_pointer == 93 && y_pointer == 75)
||(x_pointer == 94 && y_pointer == 75)
||(x_pointer == 95 && y_pointer == 75)
||(x_pointer == 96 && y_pointer == 75)
||(x_pointer == 97 && y_pointer == 75)
||(x_pointer == 98 && y_pointer == 75)
||(x_pointer == 99 && y_pointer == 75)
||(x_pointer == 100 && y_pointer == 75)
||(x_pointer == 101 && y_pointer == 75)
||(x_pointer == 102 && y_pointer == 75)
||(x_pointer == 103 && y_pointer == 75)
||(x_pointer == 104 && y_pointer == 75)
||(x_pointer == 56 && y_pointer == 76)
||(x_pointer == 57 && y_pointer == 76)
||(x_pointer == 58 && y_pointer == 76)
||(x_pointer == 59 && y_pointer == 76)
||(x_pointer == 60 && y_pointer == 76)
||(x_pointer == 61 && y_pointer == 76)
||(x_pointer == 62 && y_pointer == 76)
||(x_pointer == 63 && y_pointer == 76)
||(x_pointer == 64 && y_pointer == 76)
||(x_pointer == 65 && y_pointer == 76)
||(x_pointer == 66 && y_pointer == 76)
||(x_pointer == 67 && y_pointer == 76)
||(x_pointer == 68 && y_pointer == 76)
||(x_pointer == 69 && y_pointer == 76)
||(x_pointer == 70 && y_pointer == 76)
||(x_pointer == 71 && y_pointer == 76)
||(x_pointer == 72 && y_pointer == 76)
||(x_pointer == 73 && y_pointer == 76)
||(x_pointer == 74 && y_pointer == 76)
||(x_pointer == 75 && y_pointer == 76)
||(x_pointer == 76 && y_pointer == 76)
||(x_pointer == 77 && y_pointer == 76)
||(x_pointer == 78 && y_pointer == 76)
||(x_pointer == 79 && y_pointer == 76)
||(x_pointer == 80 && y_pointer == 76)
||(x_pointer == 81 && y_pointer == 76)
||(x_pointer == 82 && y_pointer == 76)
||(x_pointer == 83 && y_pointer == 76)
||(x_pointer == 84 && y_pointer == 76)
||(x_pointer == 85 && y_pointer == 76)
||(x_pointer == 86 && y_pointer == 76)
||(x_pointer == 87 && y_pointer == 76)
||(x_pointer == 88 && y_pointer == 76)
||(x_pointer == 89 && y_pointer == 76)
||(x_pointer == 90 && y_pointer == 76)
||(x_pointer == 91 && y_pointer == 76)
||(x_pointer == 92 && y_pointer == 76)
||(x_pointer == 93 && y_pointer == 76)
||(x_pointer == 94 && y_pointer == 76)
||(x_pointer == 95 && y_pointer == 76)
||(x_pointer == 96 && y_pointer == 76)
||(x_pointer == 97 && y_pointer == 76)
||(x_pointer == 98 && y_pointer == 76)
||(x_pointer == 99 && y_pointer == 76)
||(x_pointer == 100 && y_pointer == 76)
||(x_pointer == 101 && y_pointer == 76)
||(x_pointer == 102 && y_pointer == 76)
||(x_pointer == 103 && y_pointer == 76)
||(x_pointer == 104 && y_pointer == 76)
||(x_pointer == 56 && y_pointer == 77)
||(x_pointer == 57 && y_pointer == 77)
||(x_pointer == 58 && y_pointer == 77)
||(x_pointer == 59 && y_pointer == 77)
||(x_pointer == 60 && y_pointer == 77)
||(x_pointer == 61 && y_pointer == 77)
||(x_pointer == 62 && y_pointer == 77)
||(x_pointer == 63 && y_pointer == 77)
||(x_pointer == 64 && y_pointer == 77)
||(x_pointer == 65 && y_pointer == 77)
||(x_pointer == 66 && y_pointer == 77)
||(x_pointer == 67 && y_pointer == 77)
||(x_pointer == 68 && y_pointer == 77)
||(x_pointer == 69 && y_pointer == 77)
||(x_pointer == 70 && y_pointer == 77)
||(x_pointer == 71 && y_pointer == 77)
||(x_pointer == 72 && y_pointer == 77)
||(x_pointer == 73 && y_pointer == 77)
||(x_pointer == 74 && y_pointer == 77)
||(x_pointer == 75 && y_pointer == 77)
||(x_pointer == 76 && y_pointer == 77)
||(x_pointer == 77 && y_pointer == 77)
||(x_pointer == 78 && y_pointer == 77)
||(x_pointer == 79 && y_pointer == 77)
||(x_pointer == 80 && y_pointer == 77)
||(x_pointer == 81 && y_pointer == 77)
||(x_pointer == 82 && y_pointer == 77)
||(x_pointer == 83 && y_pointer == 77)
||(x_pointer == 84 && y_pointer == 77)
||(x_pointer == 85 && y_pointer == 77)
||(x_pointer == 86 && y_pointer == 77)
||(x_pointer == 87 && y_pointer == 77)
||(x_pointer == 88 && y_pointer == 77)
||(x_pointer == 89 && y_pointer == 77)
||(x_pointer == 90 && y_pointer == 77)
||(x_pointer == 91 && y_pointer == 77)
||(x_pointer == 92 && y_pointer == 77)
||(x_pointer == 93 && y_pointer == 77)
||(x_pointer == 94 && y_pointer == 77)
||(x_pointer == 95 && y_pointer == 77)
||(x_pointer == 96 && y_pointer == 77)
||(x_pointer == 97 && y_pointer == 77)
||(x_pointer == 98 && y_pointer == 77)
||(x_pointer == 99 && y_pointer == 77)
||(x_pointer == 100 && y_pointer == 77)
||(x_pointer == 101 && y_pointer == 77)
||(x_pointer == 102 && y_pointer == 77)
||(x_pointer == 103 && y_pointer == 77)
||(x_pointer == 104 && y_pointer == 77)
||(x_pointer == 56 && y_pointer == 78)
||(x_pointer == 57 && y_pointer == 78)
||(x_pointer == 58 && y_pointer == 78)
||(x_pointer == 59 && y_pointer == 78)
||(x_pointer == 60 && y_pointer == 78)
||(x_pointer == 61 && y_pointer == 78)
||(x_pointer == 62 && y_pointer == 78)
||(x_pointer == 63 && y_pointer == 78)
||(x_pointer == 64 && y_pointer == 78)
||(x_pointer == 65 && y_pointer == 78)
||(x_pointer == 66 && y_pointer == 78)
||(x_pointer == 67 && y_pointer == 78)
||(x_pointer == 68 && y_pointer == 78)
||(x_pointer == 69 && y_pointer == 78)
||(x_pointer == 70 && y_pointer == 78)
||(x_pointer == 71 && y_pointer == 78)
||(x_pointer == 72 && y_pointer == 78)
||(x_pointer == 73 && y_pointer == 78)
||(x_pointer == 74 && y_pointer == 78)
||(x_pointer == 75 && y_pointer == 78)
||(x_pointer == 76 && y_pointer == 78)
||(x_pointer == 77 && y_pointer == 78)
||(x_pointer == 78 && y_pointer == 78)
||(x_pointer == 79 && y_pointer == 78)
||(x_pointer == 80 && y_pointer == 78)
||(x_pointer == 81 && y_pointer == 78)
||(x_pointer == 82 && y_pointer == 78)
||(x_pointer == 83 && y_pointer == 78)
||(x_pointer == 84 && y_pointer == 78)
||(x_pointer == 85 && y_pointer == 78)
||(x_pointer == 86 && y_pointer == 78)
||(x_pointer == 87 && y_pointer == 78)
||(x_pointer == 88 && y_pointer == 78)
||(x_pointer == 89 && y_pointer == 78)
||(x_pointer == 90 && y_pointer == 78)
||(x_pointer == 91 && y_pointer == 78)
||(x_pointer == 92 && y_pointer == 78)
||(x_pointer == 93 && y_pointer == 78)
||(x_pointer == 94 && y_pointer == 78)
||(x_pointer == 95 && y_pointer == 78)
||(x_pointer == 96 && y_pointer == 78)
||(x_pointer == 97 && y_pointer == 78)
||(x_pointer == 98 && y_pointer == 78)
||(x_pointer == 99 && y_pointer == 78)
||(x_pointer == 100 && y_pointer == 78)
||(x_pointer == 101 && y_pointer == 78)
||(x_pointer == 102 && y_pointer == 78)
||(x_pointer == 103 && y_pointer == 78)
||(x_pointer == 104 && y_pointer == 78)
||(x_pointer == 56 && y_pointer == 79)
||(x_pointer == 57 && y_pointer == 79)
||(x_pointer == 58 && y_pointer == 79)
||(x_pointer == 59 && y_pointer == 79)
||(x_pointer == 60 && y_pointer == 79)
||(x_pointer == 61 && y_pointer == 79)
||(x_pointer == 62 && y_pointer == 79)
||(x_pointer == 63 && y_pointer == 79)
||(x_pointer == 64 && y_pointer == 79)
||(x_pointer == 65 && y_pointer == 79)
||(x_pointer == 66 && y_pointer == 79)
||(x_pointer == 67 && y_pointer == 79)
||(x_pointer == 68 && y_pointer == 79)
||(x_pointer == 69 && y_pointer == 79)
||(x_pointer == 70 && y_pointer == 79)
||(x_pointer == 71 && y_pointer == 79)
||(x_pointer == 72 && y_pointer == 79)
||(x_pointer == 73 && y_pointer == 79)
||(x_pointer == 74 && y_pointer == 79)
||(x_pointer == 75 && y_pointer == 79)
||(x_pointer == 76 && y_pointer == 79)
||(x_pointer == 77 && y_pointer == 79)
||(x_pointer == 78 && y_pointer == 79)
||(x_pointer == 79 && y_pointer == 79)
||(x_pointer == 80 && y_pointer == 79)
||(x_pointer == 81 && y_pointer == 79)
||(x_pointer == 82 && y_pointer == 79)
||(x_pointer == 83 && y_pointer == 79)
||(x_pointer == 84 && y_pointer == 79)
||(x_pointer == 85 && y_pointer == 79)
||(x_pointer == 86 && y_pointer == 79)
||(x_pointer == 87 && y_pointer == 79)
||(x_pointer == 88 && y_pointer == 79)
||(x_pointer == 89 && y_pointer == 79)
||(x_pointer == 90 && y_pointer == 79)
||(x_pointer == 91 && y_pointer == 79)
||(x_pointer == 92 && y_pointer == 79)
||(x_pointer == 93 && y_pointer == 79)
||(x_pointer == 94 && y_pointer == 79)
||(x_pointer == 95 && y_pointer == 79)
||(x_pointer == 96 && y_pointer == 79)
||(x_pointer == 97 && y_pointer == 79)
||(x_pointer == 98 && y_pointer == 79)
||(x_pointer == 99 && y_pointer == 79)
||(x_pointer == 100 && y_pointer == 79)
||(x_pointer == 101 && y_pointer == 79)
||(x_pointer == 102 && y_pointer == 79)
||(x_pointer == 103 && y_pointer == 79)
||(x_pointer == 104 && y_pointer == 79)
||(x_pointer == 56 && y_pointer == 80)
||(x_pointer == 57 && y_pointer == 80)
||(x_pointer == 58 && y_pointer == 80)
||(x_pointer == 59 && y_pointer == 80)
||(x_pointer == 60 && y_pointer == 80)
||(x_pointer == 61 && y_pointer == 80)
||(x_pointer == 62 && y_pointer == 80)
||(x_pointer == 63 && y_pointer == 80)
||(x_pointer == 64 && y_pointer == 80)
||(x_pointer == 65 && y_pointer == 80)
||(x_pointer == 66 && y_pointer == 80)
||(x_pointer == 67 && y_pointer == 80)
||(x_pointer == 68 && y_pointer == 80)
||(x_pointer == 69 && y_pointer == 80)
||(x_pointer == 70 && y_pointer == 80)
||(x_pointer == 71 && y_pointer == 80)
||(x_pointer == 72 && y_pointer == 80)
||(x_pointer == 73 && y_pointer == 80)
||(x_pointer == 74 && y_pointer == 80)
||(x_pointer == 75 && y_pointer == 80)
||(x_pointer == 76 && y_pointer == 80)
||(x_pointer == 77 && y_pointer == 80)
||(x_pointer == 78 && y_pointer == 80)
||(x_pointer == 79 && y_pointer == 80)
||(x_pointer == 80 && y_pointer == 80)
||(x_pointer == 81 && y_pointer == 80)
||(x_pointer == 82 && y_pointer == 80)
||(x_pointer == 83 && y_pointer == 80)
||(x_pointer == 84 && y_pointer == 80)
||(x_pointer == 85 && y_pointer == 80)
||(x_pointer == 86 && y_pointer == 80)
||(x_pointer == 87 && y_pointer == 80)
||(x_pointer == 88 && y_pointer == 80)
||(x_pointer == 89 && y_pointer == 80)
||(x_pointer == 90 && y_pointer == 80)
||(x_pointer == 91 && y_pointer == 80)
||(x_pointer == 92 && y_pointer == 80)
||(x_pointer == 93 && y_pointer == 80)
||(x_pointer == 94 && y_pointer == 80)
||(x_pointer == 95 && y_pointer == 80)
||(x_pointer == 96 && y_pointer == 80)
||(x_pointer == 97 && y_pointer == 80)
||(x_pointer == 98 && y_pointer == 80)
||(x_pointer == 99 && y_pointer == 80)
||(x_pointer == 100 && y_pointer == 80)
||(x_pointer == 101 && y_pointer == 80)
||(x_pointer == 102 && y_pointer == 80)
||(x_pointer == 103 && y_pointer == 80)
||(x_pointer == 104 && y_pointer == 80)
||(x_pointer == 56 && y_pointer == 81)
||(x_pointer == 57 && y_pointer == 81)
||(x_pointer == 58 && y_pointer == 81)
||(x_pointer == 59 && y_pointer == 81)
||(x_pointer == 60 && y_pointer == 81)
||(x_pointer == 61 && y_pointer == 81)
||(x_pointer == 62 && y_pointer == 81)
||(x_pointer == 63 && y_pointer == 81)
||(x_pointer == 64 && y_pointer == 81)
||(x_pointer == 65 && y_pointer == 81)
||(x_pointer == 66 && y_pointer == 81)
||(x_pointer == 67 && y_pointer == 81)
||(x_pointer == 68 && y_pointer == 81)
||(x_pointer == 69 && y_pointer == 81)
||(x_pointer == 70 && y_pointer == 81)
||(x_pointer == 71 && y_pointer == 81)
||(x_pointer == 72 && y_pointer == 81)
||(x_pointer == 73 && y_pointer == 81)
||(x_pointer == 74 && y_pointer == 81)
||(x_pointer == 75 && y_pointer == 81)
||(x_pointer == 76 && y_pointer == 81)
||(x_pointer == 77 && y_pointer == 81)
||(x_pointer == 78 && y_pointer == 81)
||(x_pointer == 79 && y_pointer == 81)
||(x_pointer == 80 && y_pointer == 81)
||(x_pointer == 81 && y_pointer == 81)
||(x_pointer == 82 && y_pointer == 81)
||(x_pointer == 83 && y_pointer == 81)
||(x_pointer == 84 && y_pointer == 81)
||(x_pointer == 85 && y_pointer == 81)
||(x_pointer == 86 && y_pointer == 81)
||(x_pointer == 87 && y_pointer == 81)
||(x_pointer == 88 && y_pointer == 81)
||(x_pointer == 89 && y_pointer == 81)
||(x_pointer == 90 && y_pointer == 81)
||(x_pointer == 91 && y_pointer == 81)
||(x_pointer == 92 && y_pointer == 81)
||(x_pointer == 93 && y_pointer == 81)
||(x_pointer == 94 && y_pointer == 81)
||(x_pointer == 95 && y_pointer == 81)
||(x_pointer == 96 && y_pointer == 81)
||(x_pointer == 97 && y_pointer == 81)
||(x_pointer == 98 && y_pointer == 81)
||(x_pointer == 99 && y_pointer == 81)
||(x_pointer == 100 && y_pointer == 81)
||(x_pointer == 101 && y_pointer == 81)
||(x_pointer == 102 && y_pointer == 81)
||(x_pointer == 103 && y_pointer == 81)
||(x_pointer == 104 && y_pointer == 81)
||(x_pointer == 56 && y_pointer == 82)
||(x_pointer == 57 && y_pointer == 82)
||(x_pointer == 58 && y_pointer == 82)
||(x_pointer == 59 && y_pointer == 82)
||(x_pointer == 60 && y_pointer == 82)
||(x_pointer == 61 && y_pointer == 82)
||(x_pointer == 62 && y_pointer == 82)
||(x_pointer == 63 && y_pointer == 82)
||(x_pointer == 64 && y_pointer == 82)
||(x_pointer == 65 && y_pointer == 82)
||(x_pointer == 66 && y_pointer == 82)
||(x_pointer == 67 && y_pointer == 82)
||(x_pointer == 68 && y_pointer == 82)
||(x_pointer == 69 && y_pointer == 82)
||(x_pointer == 70 && y_pointer == 82)
||(x_pointer == 71 && y_pointer == 82)
||(x_pointer == 72 && y_pointer == 82)
||(x_pointer == 73 && y_pointer == 82)
||(x_pointer == 74 && y_pointer == 82)
||(x_pointer == 75 && y_pointer == 82)
||(x_pointer == 76 && y_pointer == 82)
||(x_pointer == 77 && y_pointer == 82)
||(x_pointer == 78 && y_pointer == 82)
||(x_pointer == 79 && y_pointer == 82)
||(x_pointer == 80 && y_pointer == 82)
||(x_pointer == 81 && y_pointer == 82)
||(x_pointer == 82 && y_pointer == 82)
||(x_pointer == 83 && y_pointer == 82)
||(x_pointer == 84 && y_pointer == 82)
||(x_pointer == 85 && y_pointer == 82)
||(x_pointer == 86 && y_pointer == 82)
||(x_pointer == 87 && y_pointer == 82)
||(x_pointer == 88 && y_pointer == 82)
||(x_pointer == 89 && y_pointer == 82)
||(x_pointer == 90 && y_pointer == 82)
||(x_pointer == 91 && y_pointer == 82)
||(x_pointer == 92 && y_pointer == 82)
||(x_pointer == 93 && y_pointer == 82)
||(x_pointer == 94 && y_pointer == 82)
||(x_pointer == 95 && y_pointer == 82)
||(x_pointer == 96 && y_pointer == 82)
||(x_pointer == 97 && y_pointer == 82)
||(x_pointer == 98 && y_pointer == 82)
||(x_pointer == 99 && y_pointer == 82)
||(x_pointer == 100 && y_pointer == 82)
||(x_pointer == 101 && y_pointer == 82)
||(x_pointer == 102 && y_pointer == 82)
||(x_pointer == 103 && y_pointer == 82)
||(x_pointer == 104 && y_pointer == 82)
||(x_pointer == 56 && y_pointer == 83)
||(x_pointer == 57 && y_pointer == 83)
||(x_pointer == 58 && y_pointer == 83)
||(x_pointer == 59 && y_pointer == 83)
||(x_pointer == 60 && y_pointer == 83)
||(x_pointer == 61 && y_pointer == 83)
||(x_pointer == 62 && y_pointer == 83)
||(x_pointer == 63 && y_pointer == 83)
||(x_pointer == 64 && y_pointer == 83)
||(x_pointer == 65 && y_pointer == 83)
||(x_pointer == 66 && y_pointer == 83)
||(x_pointer == 67 && y_pointer == 83)
||(x_pointer == 68 && y_pointer == 83)
||(x_pointer == 69 && y_pointer == 83)
||(x_pointer == 70 && y_pointer == 83)
||(x_pointer == 71 && y_pointer == 83)
||(x_pointer == 72 && y_pointer == 83)
||(x_pointer == 73 && y_pointer == 83)
||(x_pointer == 74 && y_pointer == 83)
||(x_pointer == 75 && y_pointer == 83)
||(x_pointer == 76 && y_pointer == 83)
||(x_pointer == 77 && y_pointer == 83)
||(x_pointer == 78 && y_pointer == 83)
||(x_pointer == 79 && y_pointer == 83)
||(x_pointer == 80 && y_pointer == 83)
||(x_pointer == 81 && y_pointer == 83)
||(x_pointer == 82 && y_pointer == 83)
||(x_pointer == 83 && y_pointer == 83)
||(x_pointer == 84 && y_pointer == 83)
||(x_pointer == 85 && y_pointer == 83)
||(x_pointer == 86 && y_pointer == 83)
||(x_pointer == 87 && y_pointer == 83)
||(x_pointer == 88 && y_pointer == 83)
||(x_pointer == 89 && y_pointer == 83)
||(x_pointer == 90 && y_pointer == 83)
||(x_pointer == 91 && y_pointer == 83)
||(x_pointer == 92 && y_pointer == 83)
||(x_pointer == 93 && y_pointer == 83)
||(x_pointer == 94 && y_pointer == 83)
||(x_pointer == 95 && y_pointer == 83)
||(x_pointer == 96 && y_pointer == 83)
||(x_pointer == 97 && y_pointer == 83)
||(x_pointer == 98 && y_pointer == 83)
||(x_pointer == 99 && y_pointer == 83)
||(x_pointer == 100 && y_pointer == 83)
||(x_pointer == 101 && y_pointer == 83)
||(x_pointer == 102 && y_pointer == 83)
||(x_pointer == 103 && y_pointer == 83)
||(x_pointer == 104 && y_pointer == 83)
||(x_pointer == 56 && y_pointer == 84)
||(x_pointer == 57 && y_pointer == 84)
||(x_pointer == 58 && y_pointer == 84)
||(x_pointer == 59 && y_pointer == 84)
||(x_pointer == 60 && y_pointer == 84)
||(x_pointer == 61 && y_pointer == 84)
||(x_pointer == 62 && y_pointer == 84)
||(x_pointer == 63 && y_pointer == 84)
||(x_pointer == 64 && y_pointer == 84)
||(x_pointer == 65 && y_pointer == 84)
||(x_pointer == 66 && y_pointer == 84)
||(x_pointer == 67 && y_pointer == 84)
||(x_pointer == 68 && y_pointer == 84)
||(x_pointer == 69 && y_pointer == 84)
||(x_pointer == 70 && y_pointer == 84)
||(x_pointer == 71 && y_pointer == 84)
||(x_pointer == 72 && y_pointer == 84)
||(x_pointer == 73 && y_pointer == 84)
||(x_pointer == 74 && y_pointer == 84)
||(x_pointer == 75 && y_pointer == 84)
||(x_pointer == 76 && y_pointer == 84)
||(x_pointer == 77 && y_pointer == 84)
||(x_pointer == 78 && y_pointer == 84)
||(x_pointer == 79 && y_pointer == 84)
||(x_pointer == 80 && y_pointer == 84)
||(x_pointer == 81 && y_pointer == 84)
||(x_pointer == 82 && y_pointer == 84)
||(x_pointer == 83 && y_pointer == 84)
||(x_pointer == 84 && y_pointer == 84)
||(x_pointer == 85 && y_pointer == 84)
||(x_pointer == 86 && y_pointer == 84)
||(x_pointer == 87 && y_pointer == 84)
||(x_pointer == 88 && y_pointer == 84)
||(x_pointer == 89 && y_pointer == 84)
||(x_pointer == 90 && y_pointer == 84)
||(x_pointer == 91 && y_pointer == 84)
||(x_pointer == 92 && y_pointer == 84)
||(x_pointer == 93 && y_pointer == 84)
||(x_pointer == 94 && y_pointer == 84)
||(x_pointer == 95 && y_pointer == 84)
||(x_pointer == 96 && y_pointer == 84)
||(x_pointer == 97 && y_pointer == 84)
||(x_pointer == 98 && y_pointer == 84)
||(x_pointer == 99 && y_pointer == 84)
||(x_pointer == 100 && y_pointer == 84)
||(x_pointer == 101 && y_pointer == 84)
||(x_pointer == 102 && y_pointer == 84)
||(x_pointer == 103 && y_pointer == 84)
||(x_pointer == 104 && y_pointer == 84)
||(x_pointer == 56 && y_pointer == 85)
||(x_pointer == 57 && y_pointer == 85)
||(x_pointer == 58 && y_pointer == 85)
||(x_pointer == 59 && y_pointer == 85)
||(x_pointer == 60 && y_pointer == 85)
||(x_pointer == 61 && y_pointer == 85)
||(x_pointer == 62 && y_pointer == 85)
||(x_pointer == 63 && y_pointer == 85)
||(x_pointer == 64 && y_pointer == 85)
||(x_pointer == 65 && y_pointer == 85)
||(x_pointer == 66 && y_pointer == 85)
||(x_pointer == 67 && y_pointer == 85)
||(x_pointer == 68 && y_pointer == 85)
||(x_pointer == 69 && y_pointer == 85)
||(x_pointer == 70 && y_pointer == 85)
||(x_pointer == 90 && y_pointer == 85)
||(x_pointer == 91 && y_pointer == 85)
||(x_pointer == 92 && y_pointer == 85)
||(x_pointer == 93 && y_pointer == 85)
||(x_pointer == 94 && y_pointer == 85)
||(x_pointer == 95 && y_pointer == 85)
||(x_pointer == 96 && y_pointer == 85)
||(x_pointer == 97 && y_pointer == 85)
||(x_pointer == 98 && y_pointer == 85)
||(x_pointer == 99 && y_pointer == 85)
||(x_pointer == 100 && y_pointer == 85)
||(x_pointer == 101 && y_pointer == 85)
||(x_pointer == 102 && y_pointer == 85)
||(x_pointer == 103 && y_pointer == 85)
||(x_pointer == 104 && y_pointer == 85)
||(x_pointer == 56 && y_pointer == 86)
||(x_pointer == 57 && y_pointer == 86)
||(x_pointer == 58 && y_pointer == 86)
||(x_pointer == 59 && y_pointer == 86)
||(x_pointer == 60 && y_pointer == 86)
||(x_pointer == 61 && y_pointer == 86)
||(x_pointer == 62 && y_pointer == 86)
||(x_pointer == 63 && y_pointer == 86)
||(x_pointer == 64 && y_pointer == 86)
||(x_pointer == 65 && y_pointer == 86)
||(x_pointer == 66 && y_pointer == 86)
||(x_pointer == 67 && y_pointer == 86)
||(x_pointer == 68 && y_pointer == 86)
||(x_pointer == 69 && y_pointer == 86)
||(x_pointer == 70 && y_pointer == 86)
||(x_pointer == 90 && y_pointer == 86)
||(x_pointer == 91 && y_pointer == 86)
||(x_pointer == 92 && y_pointer == 86)
||(x_pointer == 93 && y_pointer == 86)
||(x_pointer == 94 && y_pointer == 86)
||(x_pointer == 95 && y_pointer == 86)
||(x_pointer == 96 && y_pointer == 86)
||(x_pointer == 97 && y_pointer == 86)
||(x_pointer == 98 && y_pointer == 86)
||(x_pointer == 99 && y_pointer == 86)
||(x_pointer == 100 && y_pointer == 86)
||(x_pointer == 101 && y_pointer == 86)
||(x_pointer == 102 && y_pointer == 86)
||(x_pointer == 103 && y_pointer == 86)
||(x_pointer == 104 && y_pointer == 86)
||(x_pointer == 56 && y_pointer == 87)
||(x_pointer == 57 && y_pointer == 87)
||(x_pointer == 58 && y_pointer == 87)
||(x_pointer == 59 && y_pointer == 87)
||(x_pointer == 60 && y_pointer == 87)
||(x_pointer == 61 && y_pointer == 87)
||(x_pointer == 62 && y_pointer == 87)
||(x_pointer == 63 && y_pointer == 87)
||(x_pointer == 64 && y_pointer == 87)
||(x_pointer == 65 && y_pointer == 87)
||(x_pointer == 66 && y_pointer == 87)
||(x_pointer == 67 && y_pointer == 87)
||(x_pointer == 68 && y_pointer == 87)
||(x_pointer == 69 && y_pointer == 87)
||(x_pointer == 70 && y_pointer == 87)
||(x_pointer == 90 && y_pointer == 87)
||(x_pointer == 91 && y_pointer == 87)
||(x_pointer == 92 && y_pointer == 87)
||(x_pointer == 93 && y_pointer == 87)
||(x_pointer == 94 && y_pointer == 87)
||(x_pointer == 95 && y_pointer == 87)
||(x_pointer == 96 && y_pointer == 87)
||(x_pointer == 97 && y_pointer == 87)
||(x_pointer == 98 && y_pointer == 87)
||(x_pointer == 99 && y_pointer == 87)
||(x_pointer == 100 && y_pointer == 87)
||(x_pointer == 101 && y_pointer == 87)
||(x_pointer == 102 && y_pointer == 87)
||(x_pointer == 103 && y_pointer == 87)
||(x_pointer == 104 && y_pointer == 87)
||(x_pointer == 56 && y_pointer == 88)
||(x_pointer == 57 && y_pointer == 88)
||(x_pointer == 58 && y_pointer == 88)
||(x_pointer == 59 && y_pointer == 88)
||(x_pointer == 60 && y_pointer == 88)
||(x_pointer == 61 && y_pointer == 88)
||(x_pointer == 62 && y_pointer == 88)
||(x_pointer == 63 && y_pointer == 88)
||(x_pointer == 64 && y_pointer == 88)
||(x_pointer == 65 && y_pointer == 88)
||(x_pointer == 66 && y_pointer == 88)
||(x_pointer == 67 && y_pointer == 88)
||(x_pointer == 68 && y_pointer == 88)
||(x_pointer == 69 && y_pointer == 88)
||(x_pointer == 70 && y_pointer == 88)
||(x_pointer == 90 && y_pointer == 88)
||(x_pointer == 91 && y_pointer == 88)
||(x_pointer == 92 && y_pointer == 88)
||(x_pointer == 93 && y_pointer == 88)
||(x_pointer == 94 && y_pointer == 88)
||(x_pointer == 95 && y_pointer == 88)
||(x_pointer == 96 && y_pointer == 88)
||(x_pointer == 97 && y_pointer == 88)
||(x_pointer == 98 && y_pointer == 88)
||(x_pointer == 99 && y_pointer == 88)
||(x_pointer == 100 && y_pointer == 88)
||(x_pointer == 101 && y_pointer == 88)
||(x_pointer == 102 && y_pointer == 88)
||(x_pointer == 103 && y_pointer == 88)
||(x_pointer == 104 && y_pointer == 88)
||(x_pointer == 56 && y_pointer == 89)
||(x_pointer == 57 && y_pointer == 89)
||(x_pointer == 58 && y_pointer == 89)
||(x_pointer == 59 && y_pointer == 89)
||(x_pointer == 60 && y_pointer == 89)
||(x_pointer == 61 && y_pointer == 89)
||(x_pointer == 62 && y_pointer == 89)
||(x_pointer == 63 && y_pointer == 89)
||(x_pointer == 64 && y_pointer == 89)
||(x_pointer == 65 && y_pointer == 89)
||(x_pointer == 66 && y_pointer == 89)
||(x_pointer == 67 && y_pointer == 89)
||(x_pointer == 68 && y_pointer == 89)
||(x_pointer == 69 && y_pointer == 89)
||(x_pointer == 70 && y_pointer == 89)
||(x_pointer == 90 && y_pointer == 89)
||(x_pointer == 91 && y_pointer == 89)
||(x_pointer == 92 && y_pointer == 89)
||(x_pointer == 93 && y_pointer == 89)
||(x_pointer == 94 && y_pointer == 89)
||(x_pointer == 95 && y_pointer == 89)
||(x_pointer == 96 && y_pointer == 89)
||(x_pointer == 97 && y_pointer == 89)
||(x_pointer == 98 && y_pointer == 89)
||(x_pointer == 99 && y_pointer == 89)
||(x_pointer == 100 && y_pointer == 89)
||(x_pointer == 101 && y_pointer == 89)
||(x_pointer == 102 && y_pointer == 89)
||(x_pointer == 103 && y_pointer == 89)
||(x_pointer == 104 && y_pointer == 89)
||(x_pointer == 56 && y_pointer == 90)
||(x_pointer == 57 && y_pointer == 90)
||(x_pointer == 58 && y_pointer == 90)
||(x_pointer == 59 && y_pointer == 90)
||(x_pointer == 60 && y_pointer == 90)
||(x_pointer == 61 && y_pointer == 90)
||(x_pointer == 62 && y_pointer == 90)
||(x_pointer == 63 && y_pointer == 90)
||(x_pointer == 64 && y_pointer == 90)
||(x_pointer == 65 && y_pointer == 90)
||(x_pointer == 66 && y_pointer == 90)
||(x_pointer == 67 && y_pointer == 90)
||(x_pointer == 68 && y_pointer == 90)
||(x_pointer == 69 && y_pointer == 90)
||(x_pointer == 70 && y_pointer == 90)
||(x_pointer == 90 && y_pointer == 90)
||(x_pointer == 91 && y_pointer == 90)
||(x_pointer == 92 && y_pointer == 90)
||(x_pointer == 93 && y_pointer == 90)
||(x_pointer == 94 && y_pointer == 90)
||(x_pointer == 95 && y_pointer == 90)
||(x_pointer == 96 && y_pointer == 90)
||(x_pointer == 97 && y_pointer == 90)
||(x_pointer == 98 && y_pointer == 90)
||(x_pointer == 99 && y_pointer == 90)
||(x_pointer == 100 && y_pointer == 90)
||(x_pointer == 101 && y_pointer == 90)
||(x_pointer == 102 && y_pointer == 90)
||(x_pointer == 103 && y_pointer == 90)
||(x_pointer == 104 && y_pointer == 90)
||(x_pointer == 56 && y_pointer == 91)
||(x_pointer == 57 && y_pointer == 91)
||(x_pointer == 58 && y_pointer == 91)
||(x_pointer == 59 && y_pointer == 91)
||(x_pointer == 60 && y_pointer == 91)
||(x_pointer == 61 && y_pointer == 91)
||(x_pointer == 62 && y_pointer == 91)
||(x_pointer == 63 && y_pointer == 91)
||(x_pointer == 64 && y_pointer == 91)
||(x_pointer == 65 && y_pointer == 91)
||(x_pointer == 66 && y_pointer == 91)
||(x_pointer == 67 && y_pointer == 91)
||(x_pointer == 68 && y_pointer == 91)
||(x_pointer == 69 && y_pointer == 91)
||(x_pointer == 70 && y_pointer == 91)
||(x_pointer == 90 && y_pointer == 91)
||(x_pointer == 91 && y_pointer == 91)
||(x_pointer == 92 && y_pointer == 91)
||(x_pointer == 93 && y_pointer == 91)
||(x_pointer == 94 && y_pointer == 91)
||(x_pointer == 95 && y_pointer == 91)
||(x_pointer == 96 && y_pointer == 91)
||(x_pointer == 97 && y_pointer == 91)
||(x_pointer == 98 && y_pointer == 91)
||(x_pointer == 99 && y_pointer == 91)
||(x_pointer == 100 && y_pointer == 91)
||(x_pointer == 101 && y_pointer == 91)
||(x_pointer == 102 && y_pointer == 91)
||(x_pointer == 103 && y_pointer == 91)
||(x_pointer == 104 && y_pointer == 91)
||(x_pointer == 56 && y_pointer == 92)
||(x_pointer == 57 && y_pointer == 92)
||(x_pointer == 58 && y_pointer == 92)
||(x_pointer == 59 && y_pointer == 92)
||(x_pointer == 60 && y_pointer == 92)
||(x_pointer == 61 && y_pointer == 92)
||(x_pointer == 62 && y_pointer == 92)
||(x_pointer == 63 && y_pointer == 92)
||(x_pointer == 64 && y_pointer == 92)
||(x_pointer == 65 && y_pointer == 92)
||(x_pointer == 66 && y_pointer == 92)
||(x_pointer == 67 && y_pointer == 92)
||(x_pointer == 68 && y_pointer == 92)
||(x_pointer == 69 && y_pointer == 92)
||(x_pointer == 70 && y_pointer == 92)
||(x_pointer == 90 && y_pointer == 92)
||(x_pointer == 91 && y_pointer == 92)
||(x_pointer == 92 && y_pointer == 92)
||(x_pointer == 93 && y_pointer == 92)
||(x_pointer == 94 && y_pointer == 92)
||(x_pointer == 95 && y_pointer == 92)
||(x_pointer == 96 && y_pointer == 92)
||(x_pointer == 97 && y_pointer == 92)
||(x_pointer == 98 && y_pointer == 92)
||(x_pointer == 99 && y_pointer == 92)
||(x_pointer == 100 && y_pointer == 92)
||(x_pointer == 101 && y_pointer == 92)
||(x_pointer == 102 && y_pointer == 92)
||(x_pointer == 103 && y_pointer == 92)
||(x_pointer == 104 && y_pointer == 92)
||(x_pointer == 56 && y_pointer == 93)
||(x_pointer == 57 && y_pointer == 93)
||(x_pointer == 58 && y_pointer == 93)
||(x_pointer == 59 && y_pointer == 93)
||(x_pointer == 60 && y_pointer == 93)
||(x_pointer == 61 && y_pointer == 93)
||(x_pointer == 62 && y_pointer == 93)
||(x_pointer == 63 && y_pointer == 93)
||(x_pointer == 64 && y_pointer == 93)
||(x_pointer == 65 && y_pointer == 93)
||(x_pointer == 66 && y_pointer == 93)
||(x_pointer == 67 && y_pointer == 93)
||(x_pointer == 68 && y_pointer == 93)
||(x_pointer == 69 && y_pointer == 93)
||(x_pointer == 70 && y_pointer == 93)
||(x_pointer == 90 && y_pointer == 93)
||(x_pointer == 91 && y_pointer == 93)
||(x_pointer == 92 && y_pointer == 93)
||(x_pointer == 93 && y_pointer == 93)
||(x_pointer == 94 && y_pointer == 93)
||(x_pointer == 95 && y_pointer == 93)
||(x_pointer == 96 && y_pointer == 93)
||(x_pointer == 97 && y_pointer == 93)
||(x_pointer == 98 && y_pointer == 93)
||(x_pointer == 99 && y_pointer == 93)
||(x_pointer == 100 && y_pointer == 93)
||(x_pointer == 101 && y_pointer == 93)
||(x_pointer == 102 && y_pointer == 93)
||(x_pointer == 103 && y_pointer == 93)
||(x_pointer == 104 && y_pointer == 93)
||(x_pointer == 56 && y_pointer == 94)
||(x_pointer == 57 && y_pointer == 94)
||(x_pointer == 58 && y_pointer == 94)
||(x_pointer == 59 && y_pointer == 94)
||(x_pointer == 60 && y_pointer == 94)
||(x_pointer == 61 && y_pointer == 94)
||(x_pointer == 62 && y_pointer == 94)
||(x_pointer == 63 && y_pointer == 94)
||(x_pointer == 64 && y_pointer == 94)
||(x_pointer == 65 && y_pointer == 94)
||(x_pointer == 66 && y_pointer == 94)
||(x_pointer == 67 && y_pointer == 94)
||(x_pointer == 68 && y_pointer == 94)
||(x_pointer == 69 && y_pointer == 94)
||(x_pointer == 70 && y_pointer == 94)
||(x_pointer == 90 && y_pointer == 94)
||(x_pointer == 91 && y_pointer == 94)
||(x_pointer == 92 && y_pointer == 94)
||(x_pointer == 93 && y_pointer == 94)
||(x_pointer == 94 && y_pointer == 94)
||(x_pointer == 95 && y_pointer == 94)
||(x_pointer == 96 && y_pointer == 94)
||(x_pointer == 97 && y_pointer == 94)
||(x_pointer == 98 && y_pointer == 94)
||(x_pointer == 99 && y_pointer == 94)
||(x_pointer == 100 && y_pointer == 94)
||(x_pointer == 101 && y_pointer == 94)
||(x_pointer == 102 && y_pointer == 94)
||(x_pointer == 103 && y_pointer == 94)
||(x_pointer == 104 && y_pointer == 94)
||(x_pointer == 56 && y_pointer == 95)
||(x_pointer == 57 && y_pointer == 95)
||(x_pointer == 58 && y_pointer == 95)
||(x_pointer == 59 && y_pointer == 95)
||(x_pointer == 60 && y_pointer == 95)
||(x_pointer == 61 && y_pointer == 95)
||(x_pointer == 62 && y_pointer == 95)
||(x_pointer == 63 && y_pointer == 95)
||(x_pointer == 64 && y_pointer == 95)
||(x_pointer == 65 && y_pointer == 95)
||(x_pointer == 66 && y_pointer == 95)
||(x_pointer == 67 && y_pointer == 95)
||(x_pointer == 68 && y_pointer == 95)
||(x_pointer == 69 && y_pointer == 95)
||(x_pointer == 70 && y_pointer == 95)
||(x_pointer == 90 && y_pointer == 95)
||(x_pointer == 91 && y_pointer == 95)
||(x_pointer == 92 && y_pointer == 95)
||(x_pointer == 93 && y_pointer == 95)
||(x_pointer == 94 && y_pointer == 95)
||(x_pointer == 95 && y_pointer == 95)
||(x_pointer == 96 && y_pointer == 95)
||(x_pointer == 97 && y_pointer == 95)
||(x_pointer == 98 && y_pointer == 95)
||(x_pointer == 99 && y_pointer == 95)
||(x_pointer == 100 && y_pointer == 95)
||(x_pointer == 101 && y_pointer == 95)
||(x_pointer == 102 && y_pointer == 95)
||(x_pointer == 103 && y_pointer == 95)
||(x_pointer == 104 && y_pointer == 95)
||(x_pointer == 56 && y_pointer == 96)
||(x_pointer == 57 && y_pointer == 96)
||(x_pointer == 58 && y_pointer == 96)
||(x_pointer == 59 && y_pointer == 96)
||(x_pointer == 60 && y_pointer == 96)
||(x_pointer == 61 && y_pointer == 96)
||(x_pointer == 62 && y_pointer == 96)
||(x_pointer == 63 && y_pointer == 96)
||(x_pointer == 64 && y_pointer == 96)
||(x_pointer == 65 && y_pointer == 96)
||(x_pointer == 66 && y_pointer == 96)
||(x_pointer == 67 && y_pointer == 96)
||(x_pointer == 68 && y_pointer == 96)
||(x_pointer == 69 && y_pointer == 96)
||(x_pointer == 70 && y_pointer == 96)
||(x_pointer == 90 && y_pointer == 96)
||(x_pointer == 91 && y_pointer == 96)
||(x_pointer == 92 && y_pointer == 96)
||(x_pointer == 93 && y_pointer == 96)
||(x_pointer == 94 && y_pointer == 96)
||(x_pointer == 95 && y_pointer == 96)
||(x_pointer == 96 && y_pointer == 96)
||(x_pointer == 97 && y_pointer == 96)
||(x_pointer == 98 && y_pointer == 96)
||(x_pointer == 99 && y_pointer == 96)
||(x_pointer == 100 && y_pointer == 96)
||(x_pointer == 101 && y_pointer == 96)
||(x_pointer == 102 && y_pointer == 96)
||(x_pointer == 103 && y_pointer == 96)
||(x_pointer == 104 && y_pointer == 96)
||(x_pointer == 56 && y_pointer == 97)
||(x_pointer == 57 && y_pointer == 97)
||(x_pointer == 58 && y_pointer == 97)
||(x_pointer == 59 && y_pointer == 97)
||(x_pointer == 60 && y_pointer == 97)
||(x_pointer == 61 && y_pointer == 97)
||(x_pointer == 62 && y_pointer == 97)
||(x_pointer == 63 && y_pointer == 97)
||(x_pointer == 64 && y_pointer == 97)
||(x_pointer == 65 && y_pointer == 97)
||(x_pointer == 66 && y_pointer == 97)
||(x_pointer == 67 && y_pointer == 97)
||(x_pointer == 68 && y_pointer == 97)
||(x_pointer == 69 && y_pointer == 97)
||(x_pointer == 70 && y_pointer == 97)
||(x_pointer == 90 && y_pointer == 97)
||(x_pointer == 91 && y_pointer == 97)
||(x_pointer == 92 && y_pointer == 97)
||(x_pointer == 93 && y_pointer == 97)
||(x_pointer == 94 && y_pointer == 97)
||(x_pointer == 95 && y_pointer == 97)
||(x_pointer == 96 && y_pointer == 97)
||(x_pointer == 97 && y_pointer == 97)
||(x_pointer == 98 && y_pointer == 97)
||(x_pointer == 99 && y_pointer == 97)
||(x_pointer == 100 && y_pointer == 97)
||(x_pointer == 101 && y_pointer == 97)
||(x_pointer == 102 && y_pointer == 97)
||(x_pointer == 103 && y_pointer == 97)
||(x_pointer == 104 && y_pointer == 97));
	wire barrier_pixel_3 = current_level == 3 && ((x_pointer == 36 && y_pointer == 23)
||(x_pointer == 37 && y_pointer == 23)
||(x_pointer == 38 && y_pointer == 23)
||(x_pointer == 39 && y_pointer == 23)
||(x_pointer == 40 && y_pointer == 23)
||(x_pointer == 41 && y_pointer == 23)
||(x_pointer == 42 && y_pointer == 23)
||(x_pointer == 43 && y_pointer == 23)
||(x_pointer == 44 && y_pointer == 23)
||(x_pointer == 45 && y_pointer == 23)
||(x_pointer == 46 && y_pointer == 23)
||(x_pointer == 47 && y_pointer == 23)
||(x_pointer == 48 && y_pointer == 23)
||(x_pointer == 49 && y_pointer == 23)
||(x_pointer == 50 && y_pointer == 23)
||(x_pointer == 51 && y_pointer == 23)
||(x_pointer == 52 && y_pointer == 23)
||(x_pointer == 53 && y_pointer == 23)
||(x_pointer == 54 && y_pointer == 23)
||(x_pointer == 55 && y_pointer == 23)
||(x_pointer == 56 && y_pointer == 23)
||(x_pointer == 57 && y_pointer == 23)
||(x_pointer == 58 && y_pointer == 23)
||(x_pointer == 59 && y_pointer == 23)
||(x_pointer == 60 && y_pointer == 23)
||(x_pointer == 67 && y_pointer == 23)
||(x_pointer == 68 && y_pointer == 23)
||(x_pointer == 69 && y_pointer == 23)
||(x_pointer == 70 && y_pointer == 23)
||(x_pointer == 71 && y_pointer == 23)
||(x_pointer == 72 && y_pointer == 23)
||(x_pointer == 73 && y_pointer == 23)
||(x_pointer == 74 && y_pointer == 23)
||(x_pointer == 75 && y_pointer == 23)
||(x_pointer == 76 && y_pointer == 23)
||(x_pointer == 77 && y_pointer == 23)
||(x_pointer == 78 && y_pointer == 23)
||(x_pointer == 79 && y_pointer == 23)
||(x_pointer == 80 && y_pointer == 23)
||(x_pointer == 81 && y_pointer == 23)
||(x_pointer == 82 && y_pointer == 23)
||(x_pointer == 83 && y_pointer == 23)
||(x_pointer == 84 && y_pointer == 23)
||(x_pointer == 85 && y_pointer == 23)
||(x_pointer == 86 && y_pointer == 23)
||(x_pointer == 87 && y_pointer == 23)
||(x_pointer == 88 && y_pointer == 23)
||(x_pointer == 89 && y_pointer == 23)
||(x_pointer == 96 && y_pointer == 23)
||(x_pointer == 97 && y_pointer == 23)
||(x_pointer == 98 && y_pointer == 23)
||(x_pointer == 99 && y_pointer == 23)
||(x_pointer == 100 && y_pointer == 23)
||(x_pointer == 101 && y_pointer == 23)
||(x_pointer == 102 && y_pointer == 23)
||(x_pointer == 103 && y_pointer == 23)
||(x_pointer == 104 && y_pointer == 23)
||(x_pointer == 105 && y_pointer == 23)
||(x_pointer == 106 && y_pointer == 23)
||(x_pointer == 107 && y_pointer == 23)
||(x_pointer == 108 && y_pointer == 23)
||(x_pointer == 109 && y_pointer == 23)
||(x_pointer == 110 && y_pointer == 23)
||(x_pointer == 111 && y_pointer == 23)
||(x_pointer == 112 && y_pointer == 23)
||(x_pointer == 113 && y_pointer == 23)
||(x_pointer == 114 && y_pointer == 23)
||(x_pointer == 115 && y_pointer == 23)
||(x_pointer == 116 && y_pointer == 23)
||(x_pointer == 117 && y_pointer == 23)
||(x_pointer == 118 && y_pointer == 23)
||(x_pointer == 119 && y_pointer == 23)
||(x_pointer == 120 && y_pointer == 23)
||(x_pointer == 36 && y_pointer == 24)
||(x_pointer == 37 && y_pointer == 24)
||(x_pointer == 38 && y_pointer == 24)
||(x_pointer == 39 && y_pointer == 24)
||(x_pointer == 40 && y_pointer == 24)
||(x_pointer == 41 && y_pointer == 24)
||(x_pointer == 42 && y_pointer == 24)
||(x_pointer == 43 && y_pointer == 24)
||(x_pointer == 44 && y_pointer == 24)
||(x_pointer == 45 && y_pointer == 24)
||(x_pointer == 46 && y_pointer == 24)
||(x_pointer == 47 && y_pointer == 24)
||(x_pointer == 48 && y_pointer == 24)
||(x_pointer == 49 && y_pointer == 24)
||(x_pointer == 50 && y_pointer == 24)
||(x_pointer == 51 && y_pointer == 24)
||(x_pointer == 52 && y_pointer == 24)
||(x_pointer == 53 && y_pointer == 24)
||(x_pointer == 54 && y_pointer == 24)
||(x_pointer == 55 && y_pointer == 24)
||(x_pointer == 56 && y_pointer == 24)
||(x_pointer == 57 && y_pointer == 24)
||(x_pointer == 58 && y_pointer == 24)
||(x_pointer == 59 && y_pointer == 24)
||(x_pointer == 60 && y_pointer == 24)
||(x_pointer == 67 && y_pointer == 24)
||(x_pointer == 68 && y_pointer == 24)
||(x_pointer == 69 && y_pointer == 24)
||(x_pointer == 70 && y_pointer == 24)
||(x_pointer == 71 && y_pointer == 24)
||(x_pointer == 72 && y_pointer == 24)
||(x_pointer == 73 && y_pointer == 24)
||(x_pointer == 74 && y_pointer == 24)
||(x_pointer == 75 && y_pointer == 24)
||(x_pointer == 76 && y_pointer == 24)
||(x_pointer == 77 && y_pointer == 24)
||(x_pointer == 78 && y_pointer == 24)
||(x_pointer == 79 && y_pointer == 24)
||(x_pointer == 80 && y_pointer == 24)
||(x_pointer == 81 && y_pointer == 24)
||(x_pointer == 82 && y_pointer == 24)
||(x_pointer == 83 && y_pointer == 24)
||(x_pointer == 84 && y_pointer == 24)
||(x_pointer == 85 && y_pointer == 24)
||(x_pointer == 86 && y_pointer == 24)
||(x_pointer == 87 && y_pointer == 24)
||(x_pointer == 88 && y_pointer == 24)
||(x_pointer == 89 && y_pointer == 24)
||(x_pointer == 96 && y_pointer == 24)
||(x_pointer == 97 && y_pointer == 24)
||(x_pointer == 98 && y_pointer == 24)
||(x_pointer == 99 && y_pointer == 24)
||(x_pointer == 100 && y_pointer == 24)
||(x_pointer == 101 && y_pointer == 24)
||(x_pointer == 102 && y_pointer == 24)
||(x_pointer == 103 && y_pointer == 24)
||(x_pointer == 104 && y_pointer == 24)
||(x_pointer == 105 && y_pointer == 24)
||(x_pointer == 106 && y_pointer == 24)
||(x_pointer == 107 && y_pointer == 24)
||(x_pointer == 108 && y_pointer == 24)
||(x_pointer == 109 && y_pointer == 24)
||(x_pointer == 110 && y_pointer == 24)
||(x_pointer == 111 && y_pointer == 24)
||(x_pointer == 112 && y_pointer == 24)
||(x_pointer == 113 && y_pointer == 24)
||(x_pointer == 114 && y_pointer == 24)
||(x_pointer == 115 && y_pointer == 24)
||(x_pointer == 116 && y_pointer == 24)
||(x_pointer == 117 && y_pointer == 24)
||(x_pointer == 118 && y_pointer == 24)
||(x_pointer == 119 && y_pointer == 24)
||(x_pointer == 120 && y_pointer == 24)
||(x_pointer == 36 && y_pointer == 25)
||(x_pointer == 37 && y_pointer == 25)
||(x_pointer == 38 && y_pointer == 25)
||(x_pointer == 39 && y_pointer == 25)
||(x_pointer == 40 && y_pointer == 25)
||(x_pointer == 41 && y_pointer == 25)
||(x_pointer == 42 && y_pointer == 25)
||(x_pointer == 43 && y_pointer == 25)
||(x_pointer == 44 && y_pointer == 25)
||(x_pointer == 45 && y_pointer == 25)
||(x_pointer == 46 && y_pointer == 25)
||(x_pointer == 47 && y_pointer == 25)
||(x_pointer == 48 && y_pointer == 25)
||(x_pointer == 49 && y_pointer == 25)
||(x_pointer == 50 && y_pointer == 25)
||(x_pointer == 51 && y_pointer == 25)
||(x_pointer == 52 && y_pointer == 25)
||(x_pointer == 53 && y_pointer == 25)
||(x_pointer == 54 && y_pointer == 25)
||(x_pointer == 55 && y_pointer == 25)
||(x_pointer == 56 && y_pointer == 25)
||(x_pointer == 57 && y_pointer == 25)
||(x_pointer == 58 && y_pointer == 25)
||(x_pointer == 59 && y_pointer == 25)
||(x_pointer == 60 && y_pointer == 25)
||(x_pointer == 67 && y_pointer == 25)
||(x_pointer == 68 && y_pointer == 25)
||(x_pointer == 69 && y_pointer == 25)
||(x_pointer == 70 && y_pointer == 25)
||(x_pointer == 71 && y_pointer == 25)
||(x_pointer == 72 && y_pointer == 25)
||(x_pointer == 73 && y_pointer == 25)
||(x_pointer == 74 && y_pointer == 25)
||(x_pointer == 75 && y_pointer == 25)
||(x_pointer == 76 && y_pointer == 25)
||(x_pointer == 77 && y_pointer == 25)
||(x_pointer == 78 && y_pointer == 25)
||(x_pointer == 79 && y_pointer == 25)
||(x_pointer == 80 && y_pointer == 25)
||(x_pointer == 81 && y_pointer == 25)
||(x_pointer == 82 && y_pointer == 25)
||(x_pointer == 83 && y_pointer == 25)
||(x_pointer == 84 && y_pointer == 25)
||(x_pointer == 85 && y_pointer == 25)
||(x_pointer == 86 && y_pointer == 25)
||(x_pointer == 87 && y_pointer == 25)
||(x_pointer == 88 && y_pointer == 25)
||(x_pointer == 89 && y_pointer == 25)
||(x_pointer == 96 && y_pointer == 25)
||(x_pointer == 97 && y_pointer == 25)
||(x_pointer == 98 && y_pointer == 25)
||(x_pointer == 99 && y_pointer == 25)
||(x_pointer == 100 && y_pointer == 25)
||(x_pointer == 101 && y_pointer == 25)
||(x_pointer == 102 && y_pointer == 25)
||(x_pointer == 103 && y_pointer == 25)
||(x_pointer == 104 && y_pointer == 25)
||(x_pointer == 105 && y_pointer == 25)
||(x_pointer == 106 && y_pointer == 25)
||(x_pointer == 107 && y_pointer == 25)
||(x_pointer == 108 && y_pointer == 25)
||(x_pointer == 109 && y_pointer == 25)
||(x_pointer == 110 && y_pointer == 25)
||(x_pointer == 111 && y_pointer == 25)
||(x_pointer == 112 && y_pointer == 25)
||(x_pointer == 113 && y_pointer == 25)
||(x_pointer == 114 && y_pointer == 25)
||(x_pointer == 115 && y_pointer == 25)
||(x_pointer == 116 && y_pointer == 25)
||(x_pointer == 117 && y_pointer == 25)
||(x_pointer == 118 && y_pointer == 25)
||(x_pointer == 119 && y_pointer == 25)
||(x_pointer == 120 && y_pointer == 25)
||(x_pointer == 36 && y_pointer == 26)
||(x_pointer == 37 && y_pointer == 26)
||(x_pointer == 38 && y_pointer == 26)
||(x_pointer == 39 && y_pointer == 26)
||(x_pointer == 40 && y_pointer == 26)
||(x_pointer == 41 && y_pointer == 26)
||(x_pointer == 42 && y_pointer == 26)
||(x_pointer == 43 && y_pointer == 26)
||(x_pointer == 44 && y_pointer == 26)
||(x_pointer == 45 && y_pointer == 26)
||(x_pointer == 46 && y_pointer == 26)
||(x_pointer == 47 && y_pointer == 26)
||(x_pointer == 48 && y_pointer == 26)
||(x_pointer == 49 && y_pointer == 26)
||(x_pointer == 50 && y_pointer == 26)
||(x_pointer == 51 && y_pointer == 26)
||(x_pointer == 52 && y_pointer == 26)
||(x_pointer == 53 && y_pointer == 26)
||(x_pointer == 54 && y_pointer == 26)
||(x_pointer == 55 && y_pointer == 26)
||(x_pointer == 56 && y_pointer == 26)
||(x_pointer == 57 && y_pointer == 26)
||(x_pointer == 58 && y_pointer == 26)
||(x_pointer == 59 && y_pointer == 26)
||(x_pointer == 60 && y_pointer == 26)
||(x_pointer == 67 && y_pointer == 26)
||(x_pointer == 68 && y_pointer == 26)
||(x_pointer == 69 && y_pointer == 26)
||(x_pointer == 70 && y_pointer == 26)
||(x_pointer == 71 && y_pointer == 26)
||(x_pointer == 72 && y_pointer == 26)
||(x_pointer == 73 && y_pointer == 26)
||(x_pointer == 74 && y_pointer == 26)
||(x_pointer == 75 && y_pointer == 26)
||(x_pointer == 76 && y_pointer == 26)
||(x_pointer == 77 && y_pointer == 26)
||(x_pointer == 78 && y_pointer == 26)
||(x_pointer == 79 && y_pointer == 26)
||(x_pointer == 80 && y_pointer == 26)
||(x_pointer == 81 && y_pointer == 26)
||(x_pointer == 82 && y_pointer == 26)
||(x_pointer == 83 && y_pointer == 26)
||(x_pointer == 84 && y_pointer == 26)
||(x_pointer == 85 && y_pointer == 26)
||(x_pointer == 86 && y_pointer == 26)
||(x_pointer == 87 && y_pointer == 26)
||(x_pointer == 88 && y_pointer == 26)
||(x_pointer == 89 && y_pointer == 26)
||(x_pointer == 96 && y_pointer == 26)
||(x_pointer == 97 && y_pointer == 26)
||(x_pointer == 98 && y_pointer == 26)
||(x_pointer == 99 && y_pointer == 26)
||(x_pointer == 100 && y_pointer == 26)
||(x_pointer == 101 && y_pointer == 26)
||(x_pointer == 102 && y_pointer == 26)
||(x_pointer == 103 && y_pointer == 26)
||(x_pointer == 104 && y_pointer == 26)
||(x_pointer == 105 && y_pointer == 26)
||(x_pointer == 106 && y_pointer == 26)
||(x_pointer == 107 && y_pointer == 26)
||(x_pointer == 108 && y_pointer == 26)
||(x_pointer == 109 && y_pointer == 26)
||(x_pointer == 110 && y_pointer == 26)
||(x_pointer == 111 && y_pointer == 26)
||(x_pointer == 112 && y_pointer == 26)
||(x_pointer == 113 && y_pointer == 26)
||(x_pointer == 114 && y_pointer == 26)
||(x_pointer == 115 && y_pointer == 26)
||(x_pointer == 116 && y_pointer == 26)
||(x_pointer == 117 && y_pointer == 26)
||(x_pointer == 118 && y_pointer == 26)
||(x_pointer == 119 && y_pointer == 26)
||(x_pointer == 120 && y_pointer == 26)
||(x_pointer == 36 && y_pointer == 27)
||(x_pointer == 37 && y_pointer == 27)
||(x_pointer == 38 && y_pointer == 27)
||(x_pointer == 39 && y_pointer == 27)
||(x_pointer == 67 && y_pointer == 27)
||(x_pointer == 68 && y_pointer == 27)
||(x_pointer == 69 && y_pointer == 27)
||(x_pointer == 70 && y_pointer == 27)
||(x_pointer == 86 && y_pointer == 27)
||(x_pointer == 87 && y_pointer == 27)
||(x_pointer == 88 && y_pointer == 27)
||(x_pointer == 89 && y_pointer == 27)
||(x_pointer == 96 && y_pointer == 27)
||(x_pointer == 97 && y_pointer == 27)
||(x_pointer == 98 && y_pointer == 27)
||(x_pointer == 99 && y_pointer == 27)
||(x_pointer == 36 && y_pointer == 28)
||(x_pointer == 37 && y_pointer == 28)
||(x_pointer == 38 && y_pointer == 28)
||(x_pointer == 39 && y_pointer == 28)
||(x_pointer == 67 && y_pointer == 28)
||(x_pointer == 68 && y_pointer == 28)
||(x_pointer == 69 && y_pointer == 28)
||(x_pointer == 70 && y_pointer == 28)
||(x_pointer == 86 && y_pointer == 28)
||(x_pointer == 87 && y_pointer == 28)
||(x_pointer == 88 && y_pointer == 28)
||(x_pointer == 89 && y_pointer == 28)
||(x_pointer == 96 && y_pointer == 28)
||(x_pointer == 97 && y_pointer == 28)
||(x_pointer == 98 && y_pointer == 28)
||(x_pointer == 99 && y_pointer == 28)
||(x_pointer == 36 && y_pointer == 29)
||(x_pointer == 37 && y_pointer == 29)
||(x_pointer == 38 && y_pointer == 29)
||(x_pointer == 39 && y_pointer == 29)
||(x_pointer == 67 && y_pointer == 29)
||(x_pointer == 68 && y_pointer == 29)
||(x_pointer == 69 && y_pointer == 29)
||(x_pointer == 70 && y_pointer == 29)
||(x_pointer == 96 && y_pointer == 29)
||(x_pointer == 97 && y_pointer == 29)
||(x_pointer == 98 && y_pointer == 29)
||(x_pointer == 99 && y_pointer == 29)
||(x_pointer == 36 && y_pointer == 30)
||(x_pointer == 37 && y_pointer == 30)
||(x_pointer == 38 && y_pointer == 30)
||(x_pointer == 39 && y_pointer == 30)
||(x_pointer == 67 && y_pointer == 30)
||(x_pointer == 68 && y_pointer == 30)
||(x_pointer == 69 && y_pointer == 30)
||(x_pointer == 70 && y_pointer == 30)
||(x_pointer == 96 && y_pointer == 30)
||(x_pointer == 97 && y_pointer == 30)
||(x_pointer == 98 && y_pointer == 30)
||(x_pointer == 99 && y_pointer == 30)
||(x_pointer == 36 && y_pointer == 31)
||(x_pointer == 37 && y_pointer == 31)
||(x_pointer == 38 && y_pointer == 31)
||(x_pointer == 39 && y_pointer == 31)
||(x_pointer == 67 && y_pointer == 31)
||(x_pointer == 68 && y_pointer == 31)
||(x_pointer == 69 && y_pointer == 31)
||(x_pointer == 70 && y_pointer == 31)
||(x_pointer == 96 && y_pointer == 31)
||(x_pointer == 97 && y_pointer == 31)
||(x_pointer == 98 && y_pointer == 31)
||(x_pointer == 99 && y_pointer == 31)
||(x_pointer == 36 && y_pointer == 32)
||(x_pointer == 37 && y_pointer == 32)
||(x_pointer == 38 && y_pointer == 32)
||(x_pointer == 39 && y_pointer == 32)
||(x_pointer == 67 && y_pointer == 32)
||(x_pointer == 68 && y_pointer == 32)
||(x_pointer == 69 && y_pointer == 32)
||(x_pointer == 70 && y_pointer == 32)
||(x_pointer == 96 && y_pointer == 32)
||(x_pointer == 97 && y_pointer == 32)
||(x_pointer == 98 && y_pointer == 32)
||(x_pointer == 99 && y_pointer == 32)
||(x_pointer == 36 && y_pointer == 33)
||(x_pointer == 37 && y_pointer == 33)
||(x_pointer == 38 && y_pointer == 33)
||(x_pointer == 39 && y_pointer == 33)
||(x_pointer == 67 && y_pointer == 33)
||(x_pointer == 68 && y_pointer == 33)
||(x_pointer == 69 && y_pointer == 33)
||(x_pointer == 70 && y_pointer == 33)
||(x_pointer == 96 && y_pointer == 33)
||(x_pointer == 97 && y_pointer == 33)
||(x_pointer == 98 && y_pointer == 33)
||(x_pointer == 99 && y_pointer == 33)
||(x_pointer == 36 && y_pointer == 34)
||(x_pointer == 37 && y_pointer == 34)
||(x_pointer == 38 && y_pointer == 34)
||(x_pointer == 39 && y_pointer == 34)
||(x_pointer == 67 && y_pointer == 34)
||(x_pointer == 68 && y_pointer == 34)
||(x_pointer == 69 && y_pointer == 34)
||(x_pointer == 70 && y_pointer == 34)
||(x_pointer == 96 && y_pointer == 34)
||(x_pointer == 97 && y_pointer == 34)
||(x_pointer == 98 && y_pointer == 34)
||(x_pointer == 99 && y_pointer == 34)
||(x_pointer == 36 && y_pointer == 35)
||(x_pointer == 37 && y_pointer == 35)
||(x_pointer == 38 && y_pointer == 35)
||(x_pointer == 39 && y_pointer == 35)
||(x_pointer == 67 && y_pointer == 35)
||(x_pointer == 68 && y_pointer == 35)
||(x_pointer == 69 && y_pointer == 35)
||(x_pointer == 70 && y_pointer == 35)
||(x_pointer == 96 && y_pointer == 35)
||(x_pointer == 97 && y_pointer == 35)
||(x_pointer == 98 && y_pointer == 35)
||(x_pointer == 99 && y_pointer == 35)
||(x_pointer == 36 && y_pointer == 36)
||(x_pointer == 37 && y_pointer == 36)
||(x_pointer == 38 && y_pointer == 36)
||(x_pointer == 39 && y_pointer == 36)
||(x_pointer == 67 && y_pointer == 36)
||(x_pointer == 68 && y_pointer == 36)
||(x_pointer == 69 && y_pointer == 36)
||(x_pointer == 70 && y_pointer == 36)
||(x_pointer == 71 && y_pointer == 36)
||(x_pointer == 72 && y_pointer == 36)
||(x_pointer == 73 && y_pointer == 36)
||(x_pointer == 74 && y_pointer == 36)
||(x_pointer == 75 && y_pointer == 36)
||(x_pointer == 76 && y_pointer == 36)
||(x_pointer == 77 && y_pointer == 36)
||(x_pointer == 78 && y_pointer == 36)
||(x_pointer == 79 && y_pointer == 36)
||(x_pointer == 80 && y_pointer == 36)
||(x_pointer == 81 && y_pointer == 36)
||(x_pointer == 82 && y_pointer == 36)
||(x_pointer == 83 && y_pointer == 36)
||(x_pointer == 84 && y_pointer == 36)
||(x_pointer == 85 && y_pointer == 36)
||(x_pointer == 86 && y_pointer == 36)
||(x_pointer == 87 && y_pointer == 36)
||(x_pointer == 88 && y_pointer == 36)
||(x_pointer == 89 && y_pointer == 36)
||(x_pointer == 96 && y_pointer == 36)
||(x_pointer == 97 && y_pointer == 36)
||(x_pointer == 98 && y_pointer == 36)
||(x_pointer == 99 && y_pointer == 36)
||(x_pointer == 36 && y_pointer == 37)
||(x_pointer == 37 && y_pointer == 37)
||(x_pointer == 38 && y_pointer == 37)
||(x_pointer == 39 && y_pointer == 37)
||(x_pointer == 67 && y_pointer == 37)
||(x_pointer == 68 && y_pointer == 37)
||(x_pointer == 69 && y_pointer == 37)
||(x_pointer == 70 && y_pointer == 37)
||(x_pointer == 71 && y_pointer == 37)
||(x_pointer == 72 && y_pointer == 37)
||(x_pointer == 73 && y_pointer == 37)
||(x_pointer == 74 && y_pointer == 37)
||(x_pointer == 75 && y_pointer == 37)
||(x_pointer == 76 && y_pointer == 37)
||(x_pointer == 77 && y_pointer == 37)
||(x_pointer == 78 && y_pointer == 37)
||(x_pointer == 79 && y_pointer == 37)
||(x_pointer == 80 && y_pointer == 37)
||(x_pointer == 81 && y_pointer == 37)
||(x_pointer == 82 && y_pointer == 37)
||(x_pointer == 83 && y_pointer == 37)
||(x_pointer == 84 && y_pointer == 37)
||(x_pointer == 85 && y_pointer == 37)
||(x_pointer == 86 && y_pointer == 37)
||(x_pointer == 87 && y_pointer == 37)
||(x_pointer == 88 && y_pointer == 37)
||(x_pointer == 89 && y_pointer == 37)
||(x_pointer == 96 && y_pointer == 37)
||(x_pointer == 97 && y_pointer == 37)
||(x_pointer == 98 && y_pointer == 37)
||(x_pointer == 99 && y_pointer == 37)
||(x_pointer == 36 && y_pointer == 38)
||(x_pointer == 37 && y_pointer == 38)
||(x_pointer == 38 && y_pointer == 38)
||(x_pointer == 39 && y_pointer == 38)
||(x_pointer == 67 && y_pointer == 38)
||(x_pointer == 68 && y_pointer == 38)
||(x_pointer == 69 && y_pointer == 38)
||(x_pointer == 70 && y_pointer == 38)
||(x_pointer == 71 && y_pointer == 38)
||(x_pointer == 72 && y_pointer == 38)
||(x_pointer == 73 && y_pointer == 38)
||(x_pointer == 74 && y_pointer == 38)
||(x_pointer == 75 && y_pointer == 38)
||(x_pointer == 76 && y_pointer == 38)
||(x_pointer == 77 && y_pointer == 38)
||(x_pointer == 78 && y_pointer == 38)
||(x_pointer == 79 && y_pointer == 38)
||(x_pointer == 80 && y_pointer == 38)
||(x_pointer == 81 && y_pointer == 38)
||(x_pointer == 82 && y_pointer == 38)
||(x_pointer == 83 && y_pointer == 38)
||(x_pointer == 84 && y_pointer == 38)
||(x_pointer == 85 && y_pointer == 38)
||(x_pointer == 86 && y_pointer == 38)
||(x_pointer == 87 && y_pointer == 38)
||(x_pointer == 88 && y_pointer == 38)
||(x_pointer == 89 && y_pointer == 38)
||(x_pointer == 96 && y_pointer == 38)
||(x_pointer == 97 && y_pointer == 38)
||(x_pointer == 98 && y_pointer == 38)
||(x_pointer == 99 && y_pointer == 38)
||(x_pointer == 36 && y_pointer == 39)
||(x_pointer == 37 && y_pointer == 39)
||(x_pointer == 38 && y_pointer == 39)
||(x_pointer == 39 && y_pointer == 39)
||(x_pointer == 67 && y_pointer == 39)
||(x_pointer == 68 && y_pointer == 39)
||(x_pointer == 69 && y_pointer == 39)
||(x_pointer == 70 && y_pointer == 39)
||(x_pointer == 71 && y_pointer == 39)
||(x_pointer == 72 && y_pointer == 39)
||(x_pointer == 73 && y_pointer == 39)
||(x_pointer == 74 && y_pointer == 39)
||(x_pointer == 75 && y_pointer == 39)
||(x_pointer == 76 && y_pointer == 39)
||(x_pointer == 77 && y_pointer == 39)
||(x_pointer == 78 && y_pointer == 39)
||(x_pointer == 79 && y_pointer == 39)
||(x_pointer == 80 && y_pointer == 39)
||(x_pointer == 81 && y_pointer == 39)
||(x_pointer == 82 && y_pointer == 39)
||(x_pointer == 83 && y_pointer == 39)
||(x_pointer == 84 && y_pointer == 39)
||(x_pointer == 85 && y_pointer == 39)
||(x_pointer == 86 && y_pointer == 39)
||(x_pointer == 87 && y_pointer == 39)
||(x_pointer == 88 && y_pointer == 39)
||(x_pointer == 89 && y_pointer == 39)
||(x_pointer == 96 && y_pointer == 39)
||(x_pointer == 97 && y_pointer == 39)
||(x_pointer == 98 && y_pointer == 39)
||(x_pointer == 99 && y_pointer == 39)
||(x_pointer == 36 && y_pointer == 40)
||(x_pointer == 37 && y_pointer == 40)
||(x_pointer == 38 && y_pointer == 40)
||(x_pointer == 39 && y_pointer == 40)
||(x_pointer == 86 && y_pointer == 40)
||(x_pointer == 87 && y_pointer == 40)
||(x_pointer == 88 && y_pointer == 40)
||(x_pointer == 89 && y_pointer == 40)
||(x_pointer == 96 && y_pointer == 40)
||(x_pointer == 97 && y_pointer == 40)
||(x_pointer == 98 && y_pointer == 40)
||(x_pointer == 99 && y_pointer == 40)
||(x_pointer == 36 && y_pointer == 41)
||(x_pointer == 37 && y_pointer == 41)
||(x_pointer == 38 && y_pointer == 41)
||(x_pointer == 39 && y_pointer == 41)
||(x_pointer == 86 && y_pointer == 41)
||(x_pointer == 87 && y_pointer == 41)
||(x_pointer == 88 && y_pointer == 41)
||(x_pointer == 89 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 99 && y_pointer == 41)
||(x_pointer == 36 && y_pointer == 42)
||(x_pointer == 37 && y_pointer == 42)
||(x_pointer == 38 && y_pointer == 42)
||(x_pointer == 39 && y_pointer == 42)
||(x_pointer == 86 && y_pointer == 42)
||(x_pointer == 87 && y_pointer == 42)
||(x_pointer == 88 && y_pointer == 42)
||(x_pointer == 89 && y_pointer == 42)
||(x_pointer == 96 && y_pointer == 42)
||(x_pointer == 97 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 99 && y_pointer == 42)
||(x_pointer == 36 && y_pointer == 43)
||(x_pointer == 37 && y_pointer == 43)
||(x_pointer == 38 && y_pointer == 43)
||(x_pointer == 39 && y_pointer == 43)
||(x_pointer == 86 && y_pointer == 43)
||(x_pointer == 87 && y_pointer == 43)
||(x_pointer == 88 && y_pointer == 43)
||(x_pointer == 89 && y_pointer == 43)
||(x_pointer == 96 && y_pointer == 43)
||(x_pointer == 97 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 99 && y_pointer == 43)
||(x_pointer == 36 && y_pointer == 44)
||(x_pointer == 37 && y_pointer == 44)
||(x_pointer == 38 && y_pointer == 44)
||(x_pointer == 39 && y_pointer == 44)
||(x_pointer == 86 && y_pointer == 44)
||(x_pointer == 87 && y_pointer == 44)
||(x_pointer == 88 && y_pointer == 44)
||(x_pointer == 89 && y_pointer == 44)
||(x_pointer == 96 && y_pointer == 44)
||(x_pointer == 97 && y_pointer == 44)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 99 && y_pointer == 44)
||(x_pointer == 36 && y_pointer == 45)
||(x_pointer == 37 && y_pointer == 45)
||(x_pointer == 38 && y_pointer == 45)
||(x_pointer == 39 && y_pointer == 45)
||(x_pointer == 86 && y_pointer == 45)
||(x_pointer == 87 && y_pointer == 45)
||(x_pointer == 88 && y_pointer == 45)
||(x_pointer == 89 && y_pointer == 45)
||(x_pointer == 96 && y_pointer == 45)
||(x_pointer == 97 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 99 && y_pointer == 45)
||(x_pointer == 36 && y_pointer == 46)
||(x_pointer == 37 && y_pointer == 46)
||(x_pointer == 38 && y_pointer == 46)
||(x_pointer == 39 && y_pointer == 46)
||(x_pointer == 86 && y_pointer == 46)
||(x_pointer == 87 && y_pointer == 46)
||(x_pointer == 88 && y_pointer == 46)
||(x_pointer == 89 && y_pointer == 46)
||(x_pointer == 96 && y_pointer == 46)
||(x_pointer == 97 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 99 && y_pointer == 46)
||(x_pointer == 36 && y_pointer == 47)
||(x_pointer == 37 && y_pointer == 47)
||(x_pointer == 38 && y_pointer == 47)
||(x_pointer == 39 && y_pointer == 47)
||(x_pointer == 67 && y_pointer == 47)
||(x_pointer == 68 && y_pointer == 47)
||(x_pointer == 69 && y_pointer == 47)
||(x_pointer == 70 && y_pointer == 47)
||(x_pointer == 86 && y_pointer == 47)
||(x_pointer == 87 && y_pointer == 47)
||(x_pointer == 88 && y_pointer == 47)
||(x_pointer == 89 && y_pointer == 47)
||(x_pointer == 96 && y_pointer == 47)
||(x_pointer == 97 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 99 && y_pointer == 47)
||(x_pointer == 36 && y_pointer == 48)
||(x_pointer == 37 && y_pointer == 48)
||(x_pointer == 38 && y_pointer == 48)
||(x_pointer == 39 && y_pointer == 48)
||(x_pointer == 67 && y_pointer == 48)
||(x_pointer == 68 && y_pointer == 48)
||(x_pointer == 69 && y_pointer == 48)
||(x_pointer == 70 && y_pointer == 48)
||(x_pointer == 86 && y_pointer == 48)
||(x_pointer == 87 && y_pointer == 48)
||(x_pointer == 88 && y_pointer == 48)
||(x_pointer == 89 && y_pointer == 48)
||(x_pointer == 96 && y_pointer == 48)
||(x_pointer == 97 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 48)
||(x_pointer == 99 && y_pointer == 48)
||(x_pointer == 36 && y_pointer == 49)
||(x_pointer == 37 && y_pointer == 49)
||(x_pointer == 38 && y_pointer == 49)
||(x_pointer == 39 && y_pointer == 49)
||(x_pointer == 40 && y_pointer == 49)
||(x_pointer == 41 && y_pointer == 49)
||(x_pointer == 42 && y_pointer == 49)
||(x_pointer == 43 && y_pointer == 49)
||(x_pointer == 44 && y_pointer == 49)
||(x_pointer == 45 && y_pointer == 49)
||(x_pointer == 46 && y_pointer == 49)
||(x_pointer == 47 && y_pointer == 49)
||(x_pointer == 48 && y_pointer == 49)
||(x_pointer == 49 && y_pointer == 49)
||(x_pointer == 50 && y_pointer == 49)
||(x_pointer == 51 && y_pointer == 49)
||(x_pointer == 52 && y_pointer == 49)
||(x_pointer == 53 && y_pointer == 49)
||(x_pointer == 54 && y_pointer == 49)
||(x_pointer == 55 && y_pointer == 49)
||(x_pointer == 56 && y_pointer == 49)
||(x_pointer == 57 && y_pointer == 49)
||(x_pointer == 58 && y_pointer == 49)
||(x_pointer == 59 && y_pointer == 49)
||(x_pointer == 60 && y_pointer == 49)
||(x_pointer == 67 && y_pointer == 49)
||(x_pointer == 68 && y_pointer == 49)
||(x_pointer == 69 && y_pointer == 49)
||(x_pointer == 70 && y_pointer == 49)
||(x_pointer == 71 && y_pointer == 49)
||(x_pointer == 72 && y_pointer == 49)
||(x_pointer == 73 && y_pointer == 49)
||(x_pointer == 74 && y_pointer == 49)
||(x_pointer == 75 && y_pointer == 49)
||(x_pointer == 76 && y_pointer == 49)
||(x_pointer == 77 && y_pointer == 49)
||(x_pointer == 78 && y_pointer == 49)
||(x_pointer == 79 && y_pointer == 49)
||(x_pointer == 80 && y_pointer == 49)
||(x_pointer == 81 && y_pointer == 49)
||(x_pointer == 82 && y_pointer == 49)
||(x_pointer == 83 && y_pointer == 49)
||(x_pointer == 84 && y_pointer == 49)
||(x_pointer == 85 && y_pointer == 49)
||(x_pointer == 86 && y_pointer == 49)
||(x_pointer == 87 && y_pointer == 49)
||(x_pointer == 88 && y_pointer == 49)
||(x_pointer == 89 && y_pointer == 49)
||(x_pointer == 96 && y_pointer == 49)
||(x_pointer == 97 && y_pointer == 49)
||(x_pointer == 98 && y_pointer == 49)
||(x_pointer == 99 && y_pointer == 49)
||(x_pointer == 100 && y_pointer == 49)
||(x_pointer == 101 && y_pointer == 49)
||(x_pointer == 102 && y_pointer == 49)
||(x_pointer == 103 && y_pointer == 49)
||(x_pointer == 104 && y_pointer == 49)
||(x_pointer == 105 && y_pointer == 49)
||(x_pointer == 106 && y_pointer == 49)
||(x_pointer == 107 && y_pointer == 49)
||(x_pointer == 108 && y_pointer == 49)
||(x_pointer == 109 && y_pointer == 49)
||(x_pointer == 110 && y_pointer == 49)
||(x_pointer == 111 && y_pointer == 49)
||(x_pointer == 112 && y_pointer == 49)
||(x_pointer == 113 && y_pointer == 49)
||(x_pointer == 114 && y_pointer == 49)
||(x_pointer == 115 && y_pointer == 49)
||(x_pointer == 116 && y_pointer == 49)
||(x_pointer == 117 && y_pointer == 49)
||(x_pointer == 118 && y_pointer == 49)
||(x_pointer == 119 && y_pointer == 49)
||(x_pointer == 120 && y_pointer == 49)
||(x_pointer == 36 && y_pointer == 50)
||(x_pointer == 37 && y_pointer == 50)
||(x_pointer == 38 && y_pointer == 50)
||(x_pointer == 39 && y_pointer == 50)
||(x_pointer == 40 && y_pointer == 50)
||(x_pointer == 41 && y_pointer == 50)
||(x_pointer == 42 && y_pointer == 50)
||(x_pointer == 43 && y_pointer == 50)
||(x_pointer == 44 && y_pointer == 50)
||(x_pointer == 45 && y_pointer == 50)
||(x_pointer == 46 && y_pointer == 50)
||(x_pointer == 47 && y_pointer == 50)
||(x_pointer == 48 && y_pointer == 50)
||(x_pointer == 49 && y_pointer == 50)
||(x_pointer == 50 && y_pointer == 50)
||(x_pointer == 51 && y_pointer == 50)
||(x_pointer == 52 && y_pointer == 50)
||(x_pointer == 53 && y_pointer == 50)
||(x_pointer == 54 && y_pointer == 50)
||(x_pointer == 55 && y_pointer == 50)
||(x_pointer == 56 && y_pointer == 50)
||(x_pointer == 57 && y_pointer == 50)
||(x_pointer == 58 && y_pointer == 50)
||(x_pointer == 59 && y_pointer == 50)
||(x_pointer == 60 && y_pointer == 50)
||(x_pointer == 67 && y_pointer == 50)
||(x_pointer == 68 && y_pointer == 50)
||(x_pointer == 69 && y_pointer == 50)
||(x_pointer == 70 && y_pointer == 50)
||(x_pointer == 71 && y_pointer == 50)
||(x_pointer == 72 && y_pointer == 50)
||(x_pointer == 73 && y_pointer == 50)
||(x_pointer == 74 && y_pointer == 50)
||(x_pointer == 75 && y_pointer == 50)
||(x_pointer == 76 && y_pointer == 50)
||(x_pointer == 77 && y_pointer == 50)
||(x_pointer == 78 && y_pointer == 50)
||(x_pointer == 79 && y_pointer == 50)
||(x_pointer == 80 && y_pointer == 50)
||(x_pointer == 81 && y_pointer == 50)
||(x_pointer == 82 && y_pointer == 50)
||(x_pointer == 83 && y_pointer == 50)
||(x_pointer == 84 && y_pointer == 50)
||(x_pointer == 85 && y_pointer == 50)
||(x_pointer == 86 && y_pointer == 50)
||(x_pointer == 87 && y_pointer == 50)
||(x_pointer == 88 && y_pointer == 50)
||(x_pointer == 89 && y_pointer == 50)
||(x_pointer == 96 && y_pointer == 50)
||(x_pointer == 97 && y_pointer == 50)
||(x_pointer == 98 && y_pointer == 50)
||(x_pointer == 99 && y_pointer == 50)
||(x_pointer == 100 && y_pointer == 50)
||(x_pointer == 101 && y_pointer == 50)
||(x_pointer == 102 && y_pointer == 50)
||(x_pointer == 103 && y_pointer == 50)
||(x_pointer == 104 && y_pointer == 50)
||(x_pointer == 105 && y_pointer == 50)
||(x_pointer == 106 && y_pointer == 50)
||(x_pointer == 107 && y_pointer == 50)
||(x_pointer == 108 && y_pointer == 50)
||(x_pointer == 109 && y_pointer == 50)
||(x_pointer == 110 && y_pointer == 50)
||(x_pointer == 111 && y_pointer == 50)
||(x_pointer == 112 && y_pointer == 50)
||(x_pointer == 113 && y_pointer == 50)
||(x_pointer == 114 && y_pointer == 50)
||(x_pointer == 115 && y_pointer == 50)
||(x_pointer == 116 && y_pointer == 50)
||(x_pointer == 117 && y_pointer == 50)
||(x_pointer == 118 && y_pointer == 50)
||(x_pointer == 119 && y_pointer == 50)
||(x_pointer == 120 && y_pointer == 50)
||(x_pointer == 36 && y_pointer == 51)
||(x_pointer == 37 && y_pointer == 51)
||(x_pointer == 38 && y_pointer == 51)
||(x_pointer == 39 && y_pointer == 51)
||(x_pointer == 40 && y_pointer == 51)
||(x_pointer == 41 && y_pointer == 51)
||(x_pointer == 42 && y_pointer == 51)
||(x_pointer == 43 && y_pointer == 51)
||(x_pointer == 44 && y_pointer == 51)
||(x_pointer == 45 && y_pointer == 51)
||(x_pointer == 46 && y_pointer == 51)
||(x_pointer == 47 && y_pointer == 51)
||(x_pointer == 48 && y_pointer == 51)
||(x_pointer == 49 && y_pointer == 51)
||(x_pointer == 50 && y_pointer == 51)
||(x_pointer == 51 && y_pointer == 51)
||(x_pointer == 52 && y_pointer == 51)
||(x_pointer == 53 && y_pointer == 51)
||(x_pointer == 54 && y_pointer == 51)
||(x_pointer == 55 && y_pointer == 51)
||(x_pointer == 56 && y_pointer == 51)
||(x_pointer == 57 && y_pointer == 51)
||(x_pointer == 58 && y_pointer == 51)
||(x_pointer == 59 && y_pointer == 51)
||(x_pointer == 60 && y_pointer == 51)
||(x_pointer == 67 && y_pointer == 51)
||(x_pointer == 68 && y_pointer == 51)
||(x_pointer == 69 && y_pointer == 51)
||(x_pointer == 70 && y_pointer == 51)
||(x_pointer == 71 && y_pointer == 51)
||(x_pointer == 72 && y_pointer == 51)
||(x_pointer == 73 && y_pointer == 51)
||(x_pointer == 74 && y_pointer == 51)
||(x_pointer == 75 && y_pointer == 51)
||(x_pointer == 76 && y_pointer == 51)
||(x_pointer == 77 && y_pointer == 51)
||(x_pointer == 78 && y_pointer == 51)
||(x_pointer == 79 && y_pointer == 51)
||(x_pointer == 80 && y_pointer == 51)
||(x_pointer == 81 && y_pointer == 51)
||(x_pointer == 82 && y_pointer == 51)
||(x_pointer == 83 && y_pointer == 51)
||(x_pointer == 84 && y_pointer == 51)
||(x_pointer == 85 && y_pointer == 51)
||(x_pointer == 86 && y_pointer == 51)
||(x_pointer == 87 && y_pointer == 51)
||(x_pointer == 88 && y_pointer == 51)
||(x_pointer == 89 && y_pointer == 51)
||(x_pointer == 96 && y_pointer == 51)
||(x_pointer == 97 && y_pointer == 51)
||(x_pointer == 98 && y_pointer == 51)
||(x_pointer == 99 && y_pointer == 51)
||(x_pointer == 100 && y_pointer == 51)
||(x_pointer == 101 && y_pointer == 51)
||(x_pointer == 102 && y_pointer == 51)
||(x_pointer == 103 && y_pointer == 51)
||(x_pointer == 104 && y_pointer == 51)
||(x_pointer == 105 && y_pointer == 51)
||(x_pointer == 106 && y_pointer == 51)
||(x_pointer == 107 && y_pointer == 51)
||(x_pointer == 108 && y_pointer == 51)
||(x_pointer == 109 && y_pointer == 51)
||(x_pointer == 110 && y_pointer == 51)
||(x_pointer == 111 && y_pointer == 51)
||(x_pointer == 112 && y_pointer == 51)
||(x_pointer == 113 && y_pointer == 51)
||(x_pointer == 114 && y_pointer == 51)
||(x_pointer == 115 && y_pointer == 51)
||(x_pointer == 116 && y_pointer == 51)
||(x_pointer == 117 && y_pointer == 51)
||(x_pointer == 118 && y_pointer == 51)
||(x_pointer == 119 && y_pointer == 51)
||(x_pointer == 120 && y_pointer == 51)
||(x_pointer == 36 && y_pointer == 52)
||(x_pointer == 37 && y_pointer == 52)
||(x_pointer == 38 && y_pointer == 52)
||(x_pointer == 39 && y_pointer == 52)
||(x_pointer == 40 && y_pointer == 52)
||(x_pointer == 41 && y_pointer == 52)
||(x_pointer == 42 && y_pointer == 52)
||(x_pointer == 43 && y_pointer == 52)
||(x_pointer == 44 && y_pointer == 52)
||(x_pointer == 45 && y_pointer == 52)
||(x_pointer == 46 && y_pointer == 52)
||(x_pointer == 47 && y_pointer == 52)
||(x_pointer == 48 && y_pointer == 52)
||(x_pointer == 49 && y_pointer == 52)
||(x_pointer == 50 && y_pointer == 52)
||(x_pointer == 51 && y_pointer == 52)
||(x_pointer == 52 && y_pointer == 52)
||(x_pointer == 53 && y_pointer == 52)
||(x_pointer == 54 && y_pointer == 52)
||(x_pointer == 55 && y_pointer == 52)
||(x_pointer == 56 && y_pointer == 52)
||(x_pointer == 57 && y_pointer == 52)
||(x_pointer == 58 && y_pointer == 52)
||(x_pointer == 59 && y_pointer == 52)
||(x_pointer == 60 && y_pointer == 52)
||(x_pointer == 67 && y_pointer == 52)
||(x_pointer == 68 && y_pointer == 52)
||(x_pointer == 69 && y_pointer == 52)
||(x_pointer == 70 && y_pointer == 52)
||(x_pointer == 71 && y_pointer == 52)
||(x_pointer == 72 && y_pointer == 52)
||(x_pointer == 73 && y_pointer == 52)
||(x_pointer == 74 && y_pointer == 52)
||(x_pointer == 75 && y_pointer == 52)
||(x_pointer == 76 && y_pointer == 52)
||(x_pointer == 77 && y_pointer == 52)
||(x_pointer == 78 && y_pointer == 52)
||(x_pointer == 79 && y_pointer == 52)
||(x_pointer == 80 && y_pointer == 52)
||(x_pointer == 81 && y_pointer == 52)
||(x_pointer == 82 && y_pointer == 52)
||(x_pointer == 83 && y_pointer == 52)
||(x_pointer == 84 && y_pointer == 52)
||(x_pointer == 85 && y_pointer == 52)
||(x_pointer == 86 && y_pointer == 52)
||(x_pointer == 87 && y_pointer == 52)
||(x_pointer == 88 && y_pointer == 52)
||(x_pointer == 89 && y_pointer == 52)
||(x_pointer == 96 && y_pointer == 52)
||(x_pointer == 97 && y_pointer == 52)
||(x_pointer == 98 && y_pointer == 52)
||(x_pointer == 99 && y_pointer == 52)
||(x_pointer == 100 && y_pointer == 52)
||(x_pointer == 101 && y_pointer == 52)
||(x_pointer == 102 && y_pointer == 52)
||(x_pointer == 103 && y_pointer == 52)
||(x_pointer == 104 && y_pointer == 52)
||(x_pointer == 105 && y_pointer == 52)
||(x_pointer == 106 && y_pointer == 52)
||(x_pointer == 107 && y_pointer == 52)
||(x_pointer == 108 && y_pointer == 52)
||(x_pointer == 109 && y_pointer == 52)
||(x_pointer == 110 && y_pointer == 52)
||(x_pointer == 111 && y_pointer == 52)
||(x_pointer == 112 && y_pointer == 52)
||(x_pointer == 113 && y_pointer == 52)
||(x_pointer == 114 && y_pointer == 52)
||(x_pointer == 115 && y_pointer == 52)
||(x_pointer == 116 && y_pointer == 52)
||(x_pointer == 117 && y_pointer == 52)
||(x_pointer == 118 && y_pointer == 52)
||(x_pointer == 119 && y_pointer == 52)
||(x_pointer == 120 && y_pointer == 52)
||(x_pointer == 36 && y_pointer == 66)
||(x_pointer == 37 && y_pointer == 66)
||(x_pointer == 38 && y_pointer == 66)
||(x_pointer == 39 && y_pointer == 66)
||(x_pointer == 40 && y_pointer == 66)
||(x_pointer == 41 && y_pointer == 66)
||(x_pointer == 42 && y_pointer == 66)
||(x_pointer == 43 && y_pointer == 66)
||(x_pointer == 44 && y_pointer == 66)
||(x_pointer == 45 && y_pointer == 66)
||(x_pointer == 46 && y_pointer == 66)
||(x_pointer == 47 && y_pointer == 66)
||(x_pointer == 48 && y_pointer == 66)
||(x_pointer == 49 && y_pointer == 66)
||(x_pointer == 50 && y_pointer == 66)
||(x_pointer == 51 && y_pointer == 66)
||(x_pointer == 52 && y_pointer == 66)
||(x_pointer == 53 && y_pointer == 66)
||(x_pointer == 54 && y_pointer == 66)
||(x_pointer == 55 && y_pointer == 66)
||(x_pointer == 56 && y_pointer == 66)
||(x_pointer == 57 && y_pointer == 66)
||(x_pointer == 58 && y_pointer == 66)
||(x_pointer == 59 && y_pointer == 66)
||(x_pointer == 60 && y_pointer == 66)
||(x_pointer == 67 && y_pointer == 66)
||(x_pointer == 68 && y_pointer == 66)
||(x_pointer == 69 && y_pointer == 66)
||(x_pointer == 70 && y_pointer == 66)
||(x_pointer == 71 && y_pointer == 66)
||(x_pointer == 72 && y_pointer == 66)
||(x_pointer == 73 && y_pointer == 66)
||(x_pointer == 74 && y_pointer == 66)
||(x_pointer == 75 && y_pointer == 66)
||(x_pointer == 76 && y_pointer == 66)
||(x_pointer == 77 && y_pointer == 66)
||(x_pointer == 78 && y_pointer == 66)
||(x_pointer == 79 && y_pointer == 66)
||(x_pointer == 80 && y_pointer == 66)
||(x_pointer == 81 && y_pointer == 66)
||(x_pointer == 82 && y_pointer == 66)
||(x_pointer == 83 && y_pointer == 66)
||(x_pointer == 84 && y_pointer == 66)
||(x_pointer == 85 && y_pointer == 66)
||(x_pointer == 86 && y_pointer == 66)
||(x_pointer == 87 && y_pointer == 66)
||(x_pointer == 88 && y_pointer == 66)
||(x_pointer == 89 && y_pointer == 66)
||(x_pointer == 96 && y_pointer == 66)
||(x_pointer == 97 && y_pointer == 66)
||(x_pointer == 98 && y_pointer == 66)
||(x_pointer == 99 && y_pointer == 66)
||(x_pointer == 100 && y_pointer == 66)
||(x_pointer == 101 && y_pointer == 66)
||(x_pointer == 102 && y_pointer == 66)
||(x_pointer == 103 && y_pointer == 66)
||(x_pointer == 104 && y_pointer == 66)
||(x_pointer == 105 && y_pointer == 66)
||(x_pointer == 106 && y_pointer == 66)
||(x_pointer == 107 && y_pointer == 66)
||(x_pointer == 108 && y_pointer == 66)
||(x_pointer == 109 && y_pointer == 66)
||(x_pointer == 110 && y_pointer == 66)
||(x_pointer == 111 && y_pointer == 66)
||(x_pointer == 112 && y_pointer == 66)
||(x_pointer == 113 && y_pointer == 66)
||(x_pointer == 114 && y_pointer == 66)
||(x_pointer == 115 && y_pointer == 66)
||(x_pointer == 116 && y_pointer == 66)
||(x_pointer == 117 && y_pointer == 66)
||(x_pointer == 118 && y_pointer == 66)
||(x_pointer == 119 && y_pointer == 66)
||(x_pointer == 120 && y_pointer == 66)
||(x_pointer == 36 && y_pointer == 67)
||(x_pointer == 37 && y_pointer == 67)
||(x_pointer == 38 && y_pointer == 67)
||(x_pointer == 39 && y_pointer == 67)
||(x_pointer == 40 && y_pointer == 67)
||(x_pointer == 41 && y_pointer == 67)
||(x_pointer == 42 && y_pointer == 67)
||(x_pointer == 43 && y_pointer == 67)
||(x_pointer == 44 && y_pointer == 67)
||(x_pointer == 45 && y_pointer == 67)
||(x_pointer == 46 && y_pointer == 67)
||(x_pointer == 47 && y_pointer == 67)
||(x_pointer == 48 && y_pointer == 67)
||(x_pointer == 49 && y_pointer == 67)
||(x_pointer == 50 && y_pointer == 67)
||(x_pointer == 51 && y_pointer == 67)
||(x_pointer == 52 && y_pointer == 67)
||(x_pointer == 53 && y_pointer == 67)
||(x_pointer == 54 && y_pointer == 67)
||(x_pointer == 55 && y_pointer == 67)
||(x_pointer == 56 && y_pointer == 67)
||(x_pointer == 57 && y_pointer == 67)
||(x_pointer == 58 && y_pointer == 67)
||(x_pointer == 59 && y_pointer == 67)
||(x_pointer == 60 && y_pointer == 67)
||(x_pointer == 67 && y_pointer == 67)
||(x_pointer == 68 && y_pointer == 67)
||(x_pointer == 69 && y_pointer == 67)
||(x_pointer == 70 && y_pointer == 67)
||(x_pointer == 71 && y_pointer == 67)
||(x_pointer == 72 && y_pointer == 67)
||(x_pointer == 73 && y_pointer == 67)
||(x_pointer == 74 && y_pointer == 67)
||(x_pointer == 75 && y_pointer == 67)
||(x_pointer == 76 && y_pointer == 67)
||(x_pointer == 77 && y_pointer == 67)
||(x_pointer == 78 && y_pointer == 67)
||(x_pointer == 79 && y_pointer == 67)
||(x_pointer == 80 && y_pointer == 67)
||(x_pointer == 81 && y_pointer == 67)
||(x_pointer == 82 && y_pointer == 67)
||(x_pointer == 83 && y_pointer == 67)
||(x_pointer == 84 && y_pointer == 67)
||(x_pointer == 85 && y_pointer == 67)
||(x_pointer == 86 && y_pointer == 67)
||(x_pointer == 87 && y_pointer == 67)
||(x_pointer == 88 && y_pointer == 67)
||(x_pointer == 89 && y_pointer == 67)
||(x_pointer == 96 && y_pointer == 67)
||(x_pointer == 97 && y_pointer == 67)
||(x_pointer == 98 && y_pointer == 67)
||(x_pointer == 99 && y_pointer == 67)
||(x_pointer == 100 && y_pointer == 67)
||(x_pointer == 101 && y_pointer == 67)
||(x_pointer == 102 && y_pointer == 67)
||(x_pointer == 103 && y_pointer == 67)
||(x_pointer == 104 && y_pointer == 67)
||(x_pointer == 105 && y_pointer == 67)
||(x_pointer == 106 && y_pointer == 67)
||(x_pointer == 107 && y_pointer == 67)
||(x_pointer == 108 && y_pointer == 67)
||(x_pointer == 109 && y_pointer == 67)
||(x_pointer == 110 && y_pointer == 67)
||(x_pointer == 111 && y_pointer == 67)
||(x_pointer == 112 && y_pointer == 67)
||(x_pointer == 113 && y_pointer == 67)
||(x_pointer == 114 && y_pointer == 67)
||(x_pointer == 115 && y_pointer == 67)
||(x_pointer == 116 && y_pointer == 67)
||(x_pointer == 117 && y_pointer == 67)
||(x_pointer == 118 && y_pointer == 67)
||(x_pointer == 119 && y_pointer == 67)
||(x_pointer == 120 && y_pointer == 67)
||(x_pointer == 36 && y_pointer == 68)
||(x_pointer == 37 && y_pointer == 68)
||(x_pointer == 38 && y_pointer == 68)
||(x_pointer == 39 && y_pointer == 68)
||(x_pointer == 40 && y_pointer == 68)
||(x_pointer == 41 && y_pointer == 68)
||(x_pointer == 42 && y_pointer == 68)
||(x_pointer == 43 && y_pointer == 68)
||(x_pointer == 44 && y_pointer == 68)
||(x_pointer == 45 && y_pointer == 68)
||(x_pointer == 46 && y_pointer == 68)
||(x_pointer == 47 && y_pointer == 68)
||(x_pointer == 48 && y_pointer == 68)
||(x_pointer == 49 && y_pointer == 68)
||(x_pointer == 50 && y_pointer == 68)
||(x_pointer == 51 && y_pointer == 68)
||(x_pointer == 52 && y_pointer == 68)
||(x_pointer == 53 && y_pointer == 68)
||(x_pointer == 54 && y_pointer == 68)
||(x_pointer == 55 && y_pointer == 68)
||(x_pointer == 56 && y_pointer == 68)
||(x_pointer == 57 && y_pointer == 68)
||(x_pointer == 58 && y_pointer == 68)
||(x_pointer == 59 && y_pointer == 68)
||(x_pointer == 60 && y_pointer == 68)
||(x_pointer == 67 && y_pointer == 68)
||(x_pointer == 68 && y_pointer == 68)
||(x_pointer == 69 && y_pointer == 68)
||(x_pointer == 70 && y_pointer == 68)
||(x_pointer == 71 && y_pointer == 68)
||(x_pointer == 72 && y_pointer == 68)
||(x_pointer == 73 && y_pointer == 68)
||(x_pointer == 74 && y_pointer == 68)
||(x_pointer == 75 && y_pointer == 68)
||(x_pointer == 76 && y_pointer == 68)
||(x_pointer == 77 && y_pointer == 68)
||(x_pointer == 78 && y_pointer == 68)
||(x_pointer == 79 && y_pointer == 68)
||(x_pointer == 80 && y_pointer == 68)
||(x_pointer == 81 && y_pointer == 68)
||(x_pointer == 82 && y_pointer == 68)
||(x_pointer == 83 && y_pointer == 68)
||(x_pointer == 84 && y_pointer == 68)
||(x_pointer == 85 && y_pointer == 68)
||(x_pointer == 86 && y_pointer == 68)
||(x_pointer == 87 && y_pointer == 68)
||(x_pointer == 88 && y_pointer == 68)
||(x_pointer == 89 && y_pointer == 68)
||(x_pointer == 96 && y_pointer == 68)
||(x_pointer == 97 && y_pointer == 68)
||(x_pointer == 98 && y_pointer == 68)
||(x_pointer == 99 && y_pointer == 68)
||(x_pointer == 100 && y_pointer == 68)
||(x_pointer == 101 && y_pointer == 68)
||(x_pointer == 102 && y_pointer == 68)
||(x_pointer == 103 && y_pointer == 68)
||(x_pointer == 104 && y_pointer == 68)
||(x_pointer == 105 && y_pointer == 68)
||(x_pointer == 106 && y_pointer == 68)
||(x_pointer == 107 && y_pointer == 68)
||(x_pointer == 108 && y_pointer == 68)
||(x_pointer == 109 && y_pointer == 68)
||(x_pointer == 110 && y_pointer == 68)
||(x_pointer == 111 && y_pointer == 68)
||(x_pointer == 112 && y_pointer == 68)
||(x_pointer == 113 && y_pointer == 68)
||(x_pointer == 114 && y_pointer == 68)
||(x_pointer == 115 && y_pointer == 68)
||(x_pointer == 116 && y_pointer == 68)
||(x_pointer == 117 && y_pointer == 68)
||(x_pointer == 118 && y_pointer == 68)
||(x_pointer == 119 && y_pointer == 68)
||(x_pointer == 120 && y_pointer == 68)
||(x_pointer == 36 && y_pointer == 69)
||(x_pointer == 37 && y_pointer == 69)
||(x_pointer == 38 && y_pointer == 69)
||(x_pointer == 39 && y_pointer == 69)
||(x_pointer == 40 && y_pointer == 69)
||(x_pointer == 41 && y_pointer == 69)
||(x_pointer == 42 && y_pointer == 69)
||(x_pointer == 43 && y_pointer == 69)
||(x_pointer == 44 && y_pointer == 69)
||(x_pointer == 45 && y_pointer == 69)
||(x_pointer == 46 && y_pointer == 69)
||(x_pointer == 47 && y_pointer == 69)
||(x_pointer == 48 && y_pointer == 69)
||(x_pointer == 49 && y_pointer == 69)
||(x_pointer == 50 && y_pointer == 69)
||(x_pointer == 51 && y_pointer == 69)
||(x_pointer == 52 && y_pointer == 69)
||(x_pointer == 53 && y_pointer == 69)
||(x_pointer == 54 && y_pointer == 69)
||(x_pointer == 55 && y_pointer == 69)
||(x_pointer == 56 && y_pointer == 69)
||(x_pointer == 57 && y_pointer == 69)
||(x_pointer == 58 && y_pointer == 69)
||(x_pointer == 59 && y_pointer == 69)
||(x_pointer == 60 && y_pointer == 69)
||(x_pointer == 67 && y_pointer == 69)
||(x_pointer == 68 && y_pointer == 69)
||(x_pointer == 69 && y_pointer == 69)
||(x_pointer == 70 && y_pointer == 69)
||(x_pointer == 71 && y_pointer == 69)
||(x_pointer == 72 && y_pointer == 69)
||(x_pointer == 73 && y_pointer == 69)
||(x_pointer == 74 && y_pointer == 69)
||(x_pointer == 75 && y_pointer == 69)
||(x_pointer == 76 && y_pointer == 69)
||(x_pointer == 77 && y_pointer == 69)
||(x_pointer == 78 && y_pointer == 69)
||(x_pointer == 79 && y_pointer == 69)
||(x_pointer == 80 && y_pointer == 69)
||(x_pointer == 81 && y_pointer == 69)
||(x_pointer == 82 && y_pointer == 69)
||(x_pointer == 83 && y_pointer == 69)
||(x_pointer == 84 && y_pointer == 69)
||(x_pointer == 85 && y_pointer == 69)
||(x_pointer == 86 && y_pointer == 69)
||(x_pointer == 87 && y_pointer == 69)
||(x_pointer == 88 && y_pointer == 69)
||(x_pointer == 89 && y_pointer == 69)
||(x_pointer == 96 && y_pointer == 69)
||(x_pointer == 97 && y_pointer == 69)
||(x_pointer == 98 && y_pointer == 69)
||(x_pointer == 99 && y_pointer == 69)
||(x_pointer == 100 && y_pointer == 69)
||(x_pointer == 101 && y_pointer == 69)
||(x_pointer == 102 && y_pointer == 69)
||(x_pointer == 103 && y_pointer == 69)
||(x_pointer == 104 && y_pointer == 69)
||(x_pointer == 105 && y_pointer == 69)
||(x_pointer == 106 && y_pointer == 69)
||(x_pointer == 107 && y_pointer == 69)
||(x_pointer == 108 && y_pointer == 69)
||(x_pointer == 109 && y_pointer == 69)
||(x_pointer == 110 && y_pointer == 69)
||(x_pointer == 111 && y_pointer == 69)
||(x_pointer == 112 && y_pointer == 69)
||(x_pointer == 113 && y_pointer == 69)
||(x_pointer == 114 && y_pointer == 69)
||(x_pointer == 115 && y_pointer == 69)
||(x_pointer == 116 && y_pointer == 69)
||(x_pointer == 117 && y_pointer == 69)
||(x_pointer == 118 && y_pointer == 69)
||(x_pointer == 119 && y_pointer == 69)
||(x_pointer == 120 && y_pointer == 69)
||(x_pointer == 57 && y_pointer == 70)
||(x_pointer == 58 && y_pointer == 70)
||(x_pointer == 59 && y_pointer == 70)
||(x_pointer == 60 && y_pointer == 70)
||(x_pointer == 67 && y_pointer == 70)
||(x_pointer == 68 && y_pointer == 70)
||(x_pointer == 69 && y_pointer == 70)
||(x_pointer == 70 && y_pointer == 70)
||(x_pointer == 96 && y_pointer == 70)
||(x_pointer == 97 && y_pointer == 70)
||(x_pointer == 98 && y_pointer == 70)
||(x_pointer == 99 && y_pointer == 70)
||(x_pointer == 117 && y_pointer == 70)
||(x_pointer == 118 && y_pointer == 70)
||(x_pointer == 119 && y_pointer == 70)
||(x_pointer == 120 && y_pointer == 70)
||(x_pointer == 57 && y_pointer == 71)
||(x_pointer == 58 && y_pointer == 71)
||(x_pointer == 59 && y_pointer == 71)
||(x_pointer == 60 && y_pointer == 71)
||(x_pointer == 67 && y_pointer == 71)
||(x_pointer == 68 && y_pointer == 71)
||(x_pointer == 69 && y_pointer == 71)
||(x_pointer == 70 && y_pointer == 71)
||(x_pointer == 96 && y_pointer == 71)
||(x_pointer == 97 && y_pointer == 71)
||(x_pointer == 98 && y_pointer == 71)
||(x_pointer == 99 && y_pointer == 71)
||(x_pointer == 117 && y_pointer == 71)
||(x_pointer == 118 && y_pointer == 71)
||(x_pointer == 119 && y_pointer == 71)
||(x_pointer == 120 && y_pointer == 71)
||(x_pointer == 57 && y_pointer == 72)
||(x_pointer == 58 && y_pointer == 72)
||(x_pointer == 59 && y_pointer == 72)
||(x_pointer == 60 && y_pointer == 72)
||(x_pointer == 67 && y_pointer == 72)
||(x_pointer == 68 && y_pointer == 72)
||(x_pointer == 69 && y_pointer == 72)
||(x_pointer == 70 && y_pointer == 72)
||(x_pointer == 96 && y_pointer == 72)
||(x_pointer == 97 && y_pointer == 72)
||(x_pointer == 98 && y_pointer == 72)
||(x_pointer == 99 && y_pointer == 72)
||(x_pointer == 117 && y_pointer == 72)
||(x_pointer == 118 && y_pointer == 72)
||(x_pointer == 119 && y_pointer == 72)
||(x_pointer == 120 && y_pointer == 72)
||(x_pointer == 57 && y_pointer == 73)
||(x_pointer == 58 && y_pointer == 73)
||(x_pointer == 59 && y_pointer == 73)
||(x_pointer == 60 && y_pointer == 73)
||(x_pointer == 67 && y_pointer == 73)
||(x_pointer == 68 && y_pointer == 73)
||(x_pointer == 69 && y_pointer == 73)
||(x_pointer == 70 && y_pointer == 73)
||(x_pointer == 96 && y_pointer == 73)
||(x_pointer == 97 && y_pointer == 73)
||(x_pointer == 98 && y_pointer == 73)
||(x_pointer == 99 && y_pointer == 73)
||(x_pointer == 117 && y_pointer == 73)
||(x_pointer == 118 && y_pointer == 73)
||(x_pointer == 119 && y_pointer == 73)
||(x_pointer == 120 && y_pointer == 73)
||(x_pointer == 57 && y_pointer == 74)
||(x_pointer == 58 && y_pointer == 74)
||(x_pointer == 59 && y_pointer == 74)
||(x_pointer == 60 && y_pointer == 74)
||(x_pointer == 67 && y_pointer == 74)
||(x_pointer == 68 && y_pointer == 74)
||(x_pointer == 69 && y_pointer == 74)
||(x_pointer == 70 && y_pointer == 74)
||(x_pointer == 96 && y_pointer == 74)
||(x_pointer == 97 && y_pointer == 74)
||(x_pointer == 98 && y_pointer == 74)
||(x_pointer == 99 && y_pointer == 74)
||(x_pointer == 117 && y_pointer == 74)
||(x_pointer == 118 && y_pointer == 74)
||(x_pointer == 119 && y_pointer == 74)
||(x_pointer == 120 && y_pointer == 74)
||(x_pointer == 57 && y_pointer == 75)
||(x_pointer == 58 && y_pointer == 75)
||(x_pointer == 59 && y_pointer == 75)
||(x_pointer == 60 && y_pointer == 75)
||(x_pointer == 67 && y_pointer == 75)
||(x_pointer == 68 && y_pointer == 75)
||(x_pointer == 69 && y_pointer == 75)
||(x_pointer == 70 && y_pointer == 75)
||(x_pointer == 96 && y_pointer == 75)
||(x_pointer == 97 && y_pointer == 75)
||(x_pointer == 98 && y_pointer == 75)
||(x_pointer == 99 && y_pointer == 75)
||(x_pointer == 117 && y_pointer == 75)
||(x_pointer == 118 && y_pointer == 75)
||(x_pointer == 119 && y_pointer == 75)
||(x_pointer == 120 && y_pointer == 75)
||(x_pointer == 57 && y_pointer == 76)
||(x_pointer == 58 && y_pointer == 76)
||(x_pointer == 59 && y_pointer == 76)
||(x_pointer == 60 && y_pointer == 76)
||(x_pointer == 67 && y_pointer == 76)
||(x_pointer == 68 && y_pointer == 76)
||(x_pointer == 69 && y_pointer == 76)
||(x_pointer == 70 && y_pointer == 76)
||(x_pointer == 96 && y_pointer == 76)
||(x_pointer == 97 && y_pointer == 76)
||(x_pointer == 98 && y_pointer == 76)
||(x_pointer == 99 && y_pointer == 76)
||(x_pointer == 117 && y_pointer == 76)
||(x_pointer == 118 && y_pointer == 76)
||(x_pointer == 119 && y_pointer == 76)
||(x_pointer == 120 && y_pointer == 76)
||(x_pointer == 57 && y_pointer == 77)
||(x_pointer == 58 && y_pointer == 77)
||(x_pointer == 59 && y_pointer == 77)
||(x_pointer == 60 && y_pointer == 77)
||(x_pointer == 67 && y_pointer == 77)
||(x_pointer == 68 && y_pointer == 77)
||(x_pointer == 69 && y_pointer == 77)
||(x_pointer == 70 && y_pointer == 77)
||(x_pointer == 96 && y_pointer == 77)
||(x_pointer == 97 && y_pointer == 77)
||(x_pointer == 98 && y_pointer == 77)
||(x_pointer == 99 && y_pointer == 77)
||(x_pointer == 117 && y_pointer == 77)
||(x_pointer == 118 && y_pointer == 77)
||(x_pointer == 119 && y_pointer == 77)
||(x_pointer == 120 && y_pointer == 77)
||(x_pointer == 57 && y_pointer == 78)
||(x_pointer == 58 && y_pointer == 78)
||(x_pointer == 59 && y_pointer == 78)
||(x_pointer == 60 && y_pointer == 78)
||(x_pointer == 67 && y_pointer == 78)
||(x_pointer == 68 && y_pointer == 78)
||(x_pointer == 69 && y_pointer == 78)
||(x_pointer == 70 && y_pointer == 78)
||(x_pointer == 96 && y_pointer == 78)
||(x_pointer == 97 && y_pointer == 78)
||(x_pointer == 98 && y_pointer == 78)
||(x_pointer == 99 && y_pointer == 78)
||(x_pointer == 117 && y_pointer == 78)
||(x_pointer == 118 && y_pointer == 78)
||(x_pointer == 119 && y_pointer == 78)
||(x_pointer == 120 && y_pointer == 78)
||(x_pointer == 57 && y_pointer == 79)
||(x_pointer == 58 && y_pointer == 79)
||(x_pointer == 59 && y_pointer == 79)
||(x_pointer == 60 && y_pointer == 79)
||(x_pointer == 67 && y_pointer == 79)
||(x_pointer == 68 && y_pointer == 79)
||(x_pointer == 69 && y_pointer == 79)
||(x_pointer == 70 && y_pointer == 79)
||(x_pointer == 96 && y_pointer == 79)
||(x_pointer == 97 && y_pointer == 79)
||(x_pointer == 98 && y_pointer == 79)
||(x_pointer == 99 && y_pointer == 79)
||(x_pointer == 117 && y_pointer == 79)
||(x_pointer == 118 && y_pointer == 79)
||(x_pointer == 119 && y_pointer == 79)
||(x_pointer == 120 && y_pointer == 79)
||(x_pointer == 36 && y_pointer == 80)
||(x_pointer == 37 && y_pointer == 80)
||(x_pointer == 38 && y_pointer == 80)
||(x_pointer == 39 && y_pointer == 80)
||(x_pointer == 40 && y_pointer == 80)
||(x_pointer == 41 && y_pointer == 80)
||(x_pointer == 42 && y_pointer == 80)
||(x_pointer == 43 && y_pointer == 80)
||(x_pointer == 44 && y_pointer == 80)
||(x_pointer == 45 && y_pointer == 80)
||(x_pointer == 46 && y_pointer == 80)
||(x_pointer == 47 && y_pointer == 80)
||(x_pointer == 48 && y_pointer == 80)
||(x_pointer == 49 && y_pointer == 80)
||(x_pointer == 50 && y_pointer == 80)
||(x_pointer == 51 && y_pointer == 80)
||(x_pointer == 52 && y_pointer == 80)
||(x_pointer == 53 && y_pointer == 80)
||(x_pointer == 54 && y_pointer == 80)
||(x_pointer == 55 && y_pointer == 80)
||(x_pointer == 56 && y_pointer == 80)
||(x_pointer == 57 && y_pointer == 80)
||(x_pointer == 58 && y_pointer == 80)
||(x_pointer == 59 && y_pointer == 80)
||(x_pointer == 60 && y_pointer == 80)
||(x_pointer == 67 && y_pointer == 80)
||(x_pointer == 68 && y_pointer == 80)
||(x_pointer == 69 && y_pointer == 80)
||(x_pointer == 70 && y_pointer == 80)
||(x_pointer == 96 && y_pointer == 80)
||(x_pointer == 97 && y_pointer == 80)
||(x_pointer == 98 && y_pointer == 80)
||(x_pointer == 99 && y_pointer == 80)
||(x_pointer == 100 && y_pointer == 80)
||(x_pointer == 101 && y_pointer == 80)
||(x_pointer == 102 && y_pointer == 80)
||(x_pointer == 103 && y_pointer == 80)
||(x_pointer == 104 && y_pointer == 80)
||(x_pointer == 105 && y_pointer == 80)
||(x_pointer == 106 && y_pointer == 80)
||(x_pointer == 107 && y_pointer == 80)
||(x_pointer == 108 && y_pointer == 80)
||(x_pointer == 109 && y_pointer == 80)
||(x_pointer == 110 && y_pointer == 80)
||(x_pointer == 111 && y_pointer == 80)
||(x_pointer == 112 && y_pointer == 80)
||(x_pointer == 113 && y_pointer == 80)
||(x_pointer == 114 && y_pointer == 80)
||(x_pointer == 115 && y_pointer == 80)
||(x_pointer == 116 && y_pointer == 80)
||(x_pointer == 117 && y_pointer == 80)
||(x_pointer == 118 && y_pointer == 80)
||(x_pointer == 119 && y_pointer == 80)
||(x_pointer == 120 && y_pointer == 80)
||(x_pointer == 36 && y_pointer == 81)
||(x_pointer == 37 && y_pointer == 81)
||(x_pointer == 38 && y_pointer == 81)
||(x_pointer == 39 && y_pointer == 81)
||(x_pointer == 40 && y_pointer == 81)
||(x_pointer == 41 && y_pointer == 81)
||(x_pointer == 42 && y_pointer == 81)
||(x_pointer == 43 && y_pointer == 81)
||(x_pointer == 44 && y_pointer == 81)
||(x_pointer == 45 && y_pointer == 81)
||(x_pointer == 46 && y_pointer == 81)
||(x_pointer == 47 && y_pointer == 81)
||(x_pointer == 48 && y_pointer == 81)
||(x_pointer == 49 && y_pointer == 81)
||(x_pointer == 50 && y_pointer == 81)
||(x_pointer == 51 && y_pointer == 81)
||(x_pointer == 52 && y_pointer == 81)
||(x_pointer == 53 && y_pointer == 81)
||(x_pointer == 54 && y_pointer == 81)
||(x_pointer == 55 && y_pointer == 81)
||(x_pointer == 56 && y_pointer == 81)
||(x_pointer == 57 && y_pointer == 81)
||(x_pointer == 58 && y_pointer == 81)
||(x_pointer == 59 && y_pointer == 81)
||(x_pointer == 60 && y_pointer == 81)
||(x_pointer == 67 && y_pointer == 81)
||(x_pointer == 68 && y_pointer == 81)
||(x_pointer == 69 && y_pointer == 81)
||(x_pointer == 70 && y_pointer == 81)
||(x_pointer == 71 && y_pointer == 81)
||(x_pointer == 72 && y_pointer == 81)
||(x_pointer == 73 && y_pointer == 81)
||(x_pointer == 74 && y_pointer == 81)
||(x_pointer == 75 && y_pointer == 81)
||(x_pointer == 76 && y_pointer == 81)
||(x_pointer == 77 && y_pointer == 81)
||(x_pointer == 78 && y_pointer == 81)
||(x_pointer == 79 && y_pointer == 81)
||(x_pointer == 80 && y_pointer == 81)
||(x_pointer == 81 && y_pointer == 81)
||(x_pointer == 82 && y_pointer == 81)
||(x_pointer == 83 && y_pointer == 81)
||(x_pointer == 84 && y_pointer == 81)
||(x_pointer == 85 && y_pointer == 81)
||(x_pointer == 86 && y_pointer == 81)
||(x_pointer == 87 && y_pointer == 81)
||(x_pointer == 88 && y_pointer == 81)
||(x_pointer == 89 && y_pointer == 81)
||(x_pointer == 96 && y_pointer == 81)
||(x_pointer == 97 && y_pointer == 81)
||(x_pointer == 98 && y_pointer == 81)
||(x_pointer == 99 && y_pointer == 81)
||(x_pointer == 100 && y_pointer == 81)
||(x_pointer == 101 && y_pointer == 81)
||(x_pointer == 102 && y_pointer == 81)
||(x_pointer == 103 && y_pointer == 81)
||(x_pointer == 104 && y_pointer == 81)
||(x_pointer == 105 && y_pointer == 81)
||(x_pointer == 106 && y_pointer == 81)
||(x_pointer == 107 && y_pointer == 81)
||(x_pointer == 108 && y_pointer == 81)
||(x_pointer == 109 && y_pointer == 81)
||(x_pointer == 110 && y_pointer == 81)
||(x_pointer == 111 && y_pointer == 81)
||(x_pointer == 112 && y_pointer == 81)
||(x_pointer == 113 && y_pointer == 81)
||(x_pointer == 114 && y_pointer == 81)
||(x_pointer == 115 && y_pointer == 81)
||(x_pointer == 116 && y_pointer == 81)
||(x_pointer == 117 && y_pointer == 81)
||(x_pointer == 118 && y_pointer == 81)
||(x_pointer == 119 && y_pointer == 81)
||(x_pointer == 120 && y_pointer == 81)
||(x_pointer == 36 && y_pointer == 82)
||(x_pointer == 37 && y_pointer == 82)
||(x_pointer == 38 && y_pointer == 82)
||(x_pointer == 39 && y_pointer == 82)
||(x_pointer == 40 && y_pointer == 82)
||(x_pointer == 41 && y_pointer == 82)
||(x_pointer == 42 && y_pointer == 82)
||(x_pointer == 43 && y_pointer == 82)
||(x_pointer == 44 && y_pointer == 82)
||(x_pointer == 45 && y_pointer == 82)
||(x_pointer == 46 && y_pointer == 82)
||(x_pointer == 47 && y_pointer == 82)
||(x_pointer == 48 && y_pointer == 82)
||(x_pointer == 49 && y_pointer == 82)
||(x_pointer == 50 && y_pointer == 82)
||(x_pointer == 51 && y_pointer == 82)
||(x_pointer == 52 && y_pointer == 82)
||(x_pointer == 53 && y_pointer == 82)
||(x_pointer == 54 && y_pointer == 82)
||(x_pointer == 55 && y_pointer == 82)
||(x_pointer == 56 && y_pointer == 82)
||(x_pointer == 57 && y_pointer == 82)
||(x_pointer == 58 && y_pointer == 82)
||(x_pointer == 59 && y_pointer == 82)
||(x_pointer == 60 && y_pointer == 82)
||(x_pointer == 67 && y_pointer == 82)
||(x_pointer == 68 && y_pointer == 82)
||(x_pointer == 69 && y_pointer == 82)
||(x_pointer == 70 && y_pointer == 82)
||(x_pointer == 71 && y_pointer == 82)
||(x_pointer == 72 && y_pointer == 82)
||(x_pointer == 73 && y_pointer == 82)
||(x_pointer == 74 && y_pointer == 82)
||(x_pointer == 75 && y_pointer == 82)
||(x_pointer == 76 && y_pointer == 82)
||(x_pointer == 77 && y_pointer == 82)
||(x_pointer == 78 && y_pointer == 82)
||(x_pointer == 79 && y_pointer == 82)
||(x_pointer == 80 && y_pointer == 82)
||(x_pointer == 81 && y_pointer == 82)
||(x_pointer == 82 && y_pointer == 82)
||(x_pointer == 83 && y_pointer == 82)
||(x_pointer == 84 && y_pointer == 82)
||(x_pointer == 85 && y_pointer == 82)
||(x_pointer == 86 && y_pointer == 82)
||(x_pointer == 87 && y_pointer == 82)
||(x_pointer == 88 && y_pointer == 82)
||(x_pointer == 89 && y_pointer == 82)
||(x_pointer == 96 && y_pointer == 82)
||(x_pointer == 97 && y_pointer == 82)
||(x_pointer == 98 && y_pointer == 82)
||(x_pointer == 99 && y_pointer == 82)
||(x_pointer == 100 && y_pointer == 82)
||(x_pointer == 101 && y_pointer == 82)
||(x_pointer == 102 && y_pointer == 82)
||(x_pointer == 103 && y_pointer == 82)
||(x_pointer == 104 && y_pointer == 82)
||(x_pointer == 105 && y_pointer == 82)
||(x_pointer == 106 && y_pointer == 82)
||(x_pointer == 107 && y_pointer == 82)
||(x_pointer == 108 && y_pointer == 82)
||(x_pointer == 109 && y_pointer == 82)
||(x_pointer == 110 && y_pointer == 82)
||(x_pointer == 111 && y_pointer == 82)
||(x_pointer == 112 && y_pointer == 82)
||(x_pointer == 113 && y_pointer == 82)
||(x_pointer == 114 && y_pointer == 82)
||(x_pointer == 115 && y_pointer == 82)
||(x_pointer == 116 && y_pointer == 82)
||(x_pointer == 117 && y_pointer == 82)
||(x_pointer == 118 && y_pointer == 82)
||(x_pointer == 119 && y_pointer == 82)
||(x_pointer == 120 && y_pointer == 82)
||(x_pointer == 36 && y_pointer == 83)
||(x_pointer == 37 && y_pointer == 83)
||(x_pointer == 38 && y_pointer == 83)
||(x_pointer == 39 && y_pointer == 83)
||(x_pointer == 40 && y_pointer == 83)
||(x_pointer == 41 && y_pointer == 83)
||(x_pointer == 42 && y_pointer == 83)
||(x_pointer == 43 && y_pointer == 83)
||(x_pointer == 44 && y_pointer == 83)
||(x_pointer == 45 && y_pointer == 83)
||(x_pointer == 46 && y_pointer == 83)
||(x_pointer == 47 && y_pointer == 83)
||(x_pointer == 48 && y_pointer == 83)
||(x_pointer == 49 && y_pointer == 83)
||(x_pointer == 50 && y_pointer == 83)
||(x_pointer == 51 && y_pointer == 83)
||(x_pointer == 52 && y_pointer == 83)
||(x_pointer == 53 && y_pointer == 83)
||(x_pointer == 54 && y_pointer == 83)
||(x_pointer == 55 && y_pointer == 83)
||(x_pointer == 56 && y_pointer == 83)
||(x_pointer == 57 && y_pointer == 83)
||(x_pointer == 58 && y_pointer == 83)
||(x_pointer == 59 && y_pointer == 83)
||(x_pointer == 60 && y_pointer == 83)
||(x_pointer == 67 && y_pointer == 83)
||(x_pointer == 68 && y_pointer == 83)
||(x_pointer == 69 && y_pointer == 83)
||(x_pointer == 70 && y_pointer == 83)
||(x_pointer == 71 && y_pointer == 83)
||(x_pointer == 72 && y_pointer == 83)
||(x_pointer == 73 && y_pointer == 83)
||(x_pointer == 74 && y_pointer == 83)
||(x_pointer == 75 && y_pointer == 83)
||(x_pointer == 76 && y_pointer == 83)
||(x_pointer == 77 && y_pointer == 83)
||(x_pointer == 78 && y_pointer == 83)
||(x_pointer == 79 && y_pointer == 83)
||(x_pointer == 80 && y_pointer == 83)
||(x_pointer == 81 && y_pointer == 83)
||(x_pointer == 82 && y_pointer == 83)
||(x_pointer == 83 && y_pointer == 83)
||(x_pointer == 84 && y_pointer == 83)
||(x_pointer == 85 && y_pointer == 83)
||(x_pointer == 86 && y_pointer == 83)
||(x_pointer == 87 && y_pointer == 83)
||(x_pointer == 88 && y_pointer == 83)
||(x_pointer == 89 && y_pointer == 83)
||(x_pointer == 96 && y_pointer == 83)
||(x_pointer == 97 && y_pointer == 83)
||(x_pointer == 98 && y_pointer == 83)
||(x_pointer == 99 && y_pointer == 83)
||(x_pointer == 100 && y_pointer == 83)
||(x_pointer == 101 && y_pointer == 83)
||(x_pointer == 102 && y_pointer == 83)
||(x_pointer == 103 && y_pointer == 83)
||(x_pointer == 104 && y_pointer == 83)
||(x_pointer == 105 && y_pointer == 83)
||(x_pointer == 106 && y_pointer == 83)
||(x_pointer == 107 && y_pointer == 83)
||(x_pointer == 108 && y_pointer == 83)
||(x_pointer == 109 && y_pointer == 83)
||(x_pointer == 110 && y_pointer == 83)
||(x_pointer == 111 && y_pointer == 83)
||(x_pointer == 112 && y_pointer == 83)
||(x_pointer == 113 && y_pointer == 83)
||(x_pointer == 114 && y_pointer == 83)
||(x_pointer == 115 && y_pointer == 83)
||(x_pointer == 116 && y_pointer == 83)
||(x_pointer == 117 && y_pointer == 83)
||(x_pointer == 118 && y_pointer == 83)
||(x_pointer == 119 && y_pointer == 83)
||(x_pointer == 120 && y_pointer == 83)
||(x_pointer == 36 && y_pointer == 84)
||(x_pointer == 37 && y_pointer == 84)
||(x_pointer == 38 && y_pointer == 84)
||(x_pointer == 39 && y_pointer == 84)
||(x_pointer == 67 && y_pointer == 84)
||(x_pointer == 68 && y_pointer == 84)
||(x_pointer == 69 && y_pointer == 84)
||(x_pointer == 70 && y_pointer == 84)
||(x_pointer == 71 && y_pointer == 84)
||(x_pointer == 72 && y_pointer == 84)
||(x_pointer == 73 && y_pointer == 84)
||(x_pointer == 74 && y_pointer == 84)
||(x_pointer == 75 && y_pointer == 84)
||(x_pointer == 76 && y_pointer == 84)
||(x_pointer == 77 && y_pointer == 84)
||(x_pointer == 78 && y_pointer == 84)
||(x_pointer == 79 && y_pointer == 84)
||(x_pointer == 80 && y_pointer == 84)
||(x_pointer == 81 && y_pointer == 84)
||(x_pointer == 82 && y_pointer == 84)
||(x_pointer == 83 && y_pointer == 84)
||(x_pointer == 84 && y_pointer == 84)
||(x_pointer == 85 && y_pointer == 84)
||(x_pointer == 86 && y_pointer == 84)
||(x_pointer == 87 && y_pointer == 84)
||(x_pointer == 88 && y_pointer == 84)
||(x_pointer == 89 && y_pointer == 84)
||(x_pointer == 96 && y_pointer == 84)
||(x_pointer == 97 && y_pointer == 84)
||(x_pointer == 98 && y_pointer == 84)
||(x_pointer == 99 && y_pointer == 84)
||(x_pointer == 100 && y_pointer == 84)
||(x_pointer == 101 && y_pointer == 84)
||(x_pointer == 102 && y_pointer == 84)
||(x_pointer == 103 && y_pointer == 84)
||(x_pointer == 104 && y_pointer == 84)
||(x_pointer == 105 && y_pointer == 84)
||(x_pointer == 106 && y_pointer == 84)
||(x_pointer == 107 && y_pointer == 84)
||(x_pointer == 108 && y_pointer == 84)
||(x_pointer == 109 && y_pointer == 84)
||(x_pointer == 110 && y_pointer == 84)
||(x_pointer == 111 && y_pointer == 84)
||(x_pointer == 112 && y_pointer == 84)
||(x_pointer == 113 && y_pointer == 84)
||(x_pointer == 114 && y_pointer == 84)
||(x_pointer == 115 && y_pointer == 84)
||(x_pointer == 116 && y_pointer == 84)
||(x_pointer == 117 && y_pointer == 84)
||(x_pointer == 118 && y_pointer == 84)
||(x_pointer == 119 && y_pointer == 84)
||(x_pointer == 120 && y_pointer == 84)
||(x_pointer == 36 && y_pointer == 85)
||(x_pointer == 37 && y_pointer == 85)
||(x_pointer == 38 && y_pointer == 85)
||(x_pointer == 39 && y_pointer == 85)
||(x_pointer == 86 && y_pointer == 85)
||(x_pointer == 87 && y_pointer == 85)
||(x_pointer == 88 && y_pointer == 85)
||(x_pointer == 89 && y_pointer == 85)
||(x_pointer == 96 && y_pointer == 85)
||(x_pointer == 97 && y_pointer == 85)
||(x_pointer == 98 && y_pointer == 85)
||(x_pointer == 99 && y_pointer == 85)
||(x_pointer == 117 && y_pointer == 85)
||(x_pointer == 118 && y_pointer == 85)
||(x_pointer == 119 && y_pointer == 85)
||(x_pointer == 120 && y_pointer == 85)
||(x_pointer == 36 && y_pointer == 86)
||(x_pointer == 37 && y_pointer == 86)
||(x_pointer == 38 && y_pointer == 86)
||(x_pointer == 39 && y_pointer == 86)
||(x_pointer == 86 && y_pointer == 86)
||(x_pointer == 87 && y_pointer == 86)
||(x_pointer == 88 && y_pointer == 86)
||(x_pointer == 89 && y_pointer == 86)
||(x_pointer == 96 && y_pointer == 86)
||(x_pointer == 97 && y_pointer == 86)
||(x_pointer == 98 && y_pointer == 86)
||(x_pointer == 99 && y_pointer == 86)
||(x_pointer == 117 && y_pointer == 86)
||(x_pointer == 118 && y_pointer == 86)
||(x_pointer == 119 && y_pointer == 86)
||(x_pointer == 120 && y_pointer == 86)
||(x_pointer == 36 && y_pointer == 87)
||(x_pointer == 37 && y_pointer == 87)
||(x_pointer == 38 && y_pointer == 87)
||(x_pointer == 39 && y_pointer == 87)
||(x_pointer == 86 && y_pointer == 87)
||(x_pointer == 87 && y_pointer == 87)
||(x_pointer == 88 && y_pointer == 87)
||(x_pointer == 89 && y_pointer == 87)
||(x_pointer == 96 && y_pointer == 87)
||(x_pointer == 97 && y_pointer == 87)
||(x_pointer == 98 && y_pointer == 87)
||(x_pointer == 99 && y_pointer == 87)
||(x_pointer == 117 && y_pointer == 87)
||(x_pointer == 118 && y_pointer == 87)
||(x_pointer == 119 && y_pointer == 87)
||(x_pointer == 120 && y_pointer == 87)
||(x_pointer == 36 && y_pointer == 88)
||(x_pointer == 37 && y_pointer == 88)
||(x_pointer == 38 && y_pointer == 88)
||(x_pointer == 39 && y_pointer == 88)
||(x_pointer == 86 && y_pointer == 88)
||(x_pointer == 87 && y_pointer == 88)
||(x_pointer == 88 && y_pointer == 88)
||(x_pointer == 89 && y_pointer == 88)
||(x_pointer == 96 && y_pointer == 88)
||(x_pointer == 97 && y_pointer == 88)
||(x_pointer == 98 && y_pointer == 88)
||(x_pointer == 99 && y_pointer == 88)
||(x_pointer == 117 && y_pointer == 88)
||(x_pointer == 118 && y_pointer == 88)
||(x_pointer == 119 && y_pointer == 88)
||(x_pointer == 120 && y_pointer == 88)
||(x_pointer == 36 && y_pointer == 89)
||(x_pointer == 37 && y_pointer == 89)
||(x_pointer == 38 && y_pointer == 89)
||(x_pointer == 39 && y_pointer == 89)
||(x_pointer == 86 && y_pointer == 89)
||(x_pointer == 87 && y_pointer == 89)
||(x_pointer == 88 && y_pointer == 89)
||(x_pointer == 89 && y_pointer == 89)
||(x_pointer == 96 && y_pointer == 89)
||(x_pointer == 97 && y_pointer == 89)
||(x_pointer == 98 && y_pointer == 89)
||(x_pointer == 99 && y_pointer == 89)
||(x_pointer == 117 && y_pointer == 89)
||(x_pointer == 118 && y_pointer == 89)
||(x_pointer == 119 && y_pointer == 89)
||(x_pointer == 120 && y_pointer == 89)
||(x_pointer == 36 && y_pointer == 90)
||(x_pointer == 37 && y_pointer == 90)
||(x_pointer == 38 && y_pointer == 90)
||(x_pointer == 39 && y_pointer == 90)
||(x_pointer == 86 && y_pointer == 90)
||(x_pointer == 87 && y_pointer == 90)
||(x_pointer == 88 && y_pointer == 90)
||(x_pointer == 89 && y_pointer == 90)
||(x_pointer == 96 && y_pointer == 90)
||(x_pointer == 97 && y_pointer == 90)
||(x_pointer == 98 && y_pointer == 90)
||(x_pointer == 99 && y_pointer == 90)
||(x_pointer == 117 && y_pointer == 90)
||(x_pointer == 118 && y_pointer == 90)
||(x_pointer == 119 && y_pointer == 90)
||(x_pointer == 120 && y_pointer == 90)
||(x_pointer == 36 && y_pointer == 91)
||(x_pointer == 37 && y_pointer == 91)
||(x_pointer == 38 && y_pointer == 91)
||(x_pointer == 39 && y_pointer == 91)
||(x_pointer == 86 && y_pointer == 91)
||(x_pointer == 87 && y_pointer == 91)
||(x_pointer == 88 && y_pointer == 91)
||(x_pointer == 89 && y_pointer == 91)
||(x_pointer == 96 && y_pointer == 91)
||(x_pointer == 97 && y_pointer == 91)
||(x_pointer == 98 && y_pointer == 91)
||(x_pointer == 99 && y_pointer == 91)
||(x_pointer == 117 && y_pointer == 91)
||(x_pointer == 118 && y_pointer == 91)
||(x_pointer == 119 && y_pointer == 91)
||(x_pointer == 120 && y_pointer == 91)
||(x_pointer == 36 && y_pointer == 92)
||(x_pointer == 37 && y_pointer == 92)
||(x_pointer == 38 && y_pointer == 92)
||(x_pointer == 39 && y_pointer == 92)
||(x_pointer == 86 && y_pointer == 92)
||(x_pointer == 87 && y_pointer == 92)
||(x_pointer == 88 && y_pointer == 92)
||(x_pointer == 89 && y_pointer == 92)
||(x_pointer == 96 && y_pointer == 92)
||(x_pointer == 97 && y_pointer == 92)
||(x_pointer == 98 && y_pointer == 92)
||(x_pointer == 99 && y_pointer == 92)
||(x_pointer == 117 && y_pointer == 92)
||(x_pointer == 118 && y_pointer == 92)
||(x_pointer == 119 && y_pointer == 92)
||(x_pointer == 120 && y_pointer == 92)
||(x_pointer == 36 && y_pointer == 93)
||(x_pointer == 37 && y_pointer == 93)
||(x_pointer == 38 && y_pointer == 93)
||(x_pointer == 39 && y_pointer == 93)
||(x_pointer == 86 && y_pointer == 93)
||(x_pointer == 87 && y_pointer == 93)
||(x_pointer == 88 && y_pointer == 93)
||(x_pointer == 89 && y_pointer == 93)
||(x_pointer == 96 && y_pointer == 93)
||(x_pointer == 97 && y_pointer == 93)
||(x_pointer == 98 && y_pointer == 93)
||(x_pointer == 99 && y_pointer == 93)
||(x_pointer == 117 && y_pointer == 93)
||(x_pointer == 118 && y_pointer == 93)
||(x_pointer == 119 && y_pointer == 93)
||(x_pointer == 120 && y_pointer == 93)
||(x_pointer == 36 && y_pointer == 94)
||(x_pointer == 37 && y_pointer == 94)
||(x_pointer == 38 && y_pointer == 94)
||(x_pointer == 39 && y_pointer == 94)
||(x_pointer == 40 && y_pointer == 94)
||(x_pointer == 41 && y_pointer == 94)
||(x_pointer == 42 && y_pointer == 94)
||(x_pointer == 43 && y_pointer == 94)
||(x_pointer == 44 && y_pointer == 94)
||(x_pointer == 45 && y_pointer == 94)
||(x_pointer == 46 && y_pointer == 94)
||(x_pointer == 47 && y_pointer == 94)
||(x_pointer == 48 && y_pointer == 94)
||(x_pointer == 49 && y_pointer == 94)
||(x_pointer == 50 && y_pointer == 94)
||(x_pointer == 51 && y_pointer == 94)
||(x_pointer == 52 && y_pointer == 94)
||(x_pointer == 53 && y_pointer == 94)
||(x_pointer == 54 && y_pointer == 94)
||(x_pointer == 55 && y_pointer == 94)
||(x_pointer == 56 && y_pointer == 94)
||(x_pointer == 57 && y_pointer == 94)
||(x_pointer == 58 && y_pointer == 94)
||(x_pointer == 59 && y_pointer == 94)
||(x_pointer == 60 && y_pointer == 94)
||(x_pointer == 67 && y_pointer == 94)
||(x_pointer == 68 && y_pointer == 94)
||(x_pointer == 69 && y_pointer == 94)
||(x_pointer == 70 && y_pointer == 94)
||(x_pointer == 71 && y_pointer == 94)
||(x_pointer == 72 && y_pointer == 94)
||(x_pointer == 73 && y_pointer == 94)
||(x_pointer == 74 && y_pointer == 94)
||(x_pointer == 75 && y_pointer == 94)
||(x_pointer == 76 && y_pointer == 94)
||(x_pointer == 77 && y_pointer == 94)
||(x_pointer == 78 && y_pointer == 94)
||(x_pointer == 79 && y_pointer == 94)
||(x_pointer == 80 && y_pointer == 94)
||(x_pointer == 81 && y_pointer == 94)
||(x_pointer == 82 && y_pointer == 94)
||(x_pointer == 83 && y_pointer == 94)
||(x_pointer == 84 && y_pointer == 94)
||(x_pointer == 85 && y_pointer == 94)
||(x_pointer == 86 && y_pointer == 94)
||(x_pointer == 87 && y_pointer == 94)
||(x_pointer == 88 && y_pointer == 94)
||(x_pointer == 89 && y_pointer == 94)
||(x_pointer == 96 && y_pointer == 94)
||(x_pointer == 97 && y_pointer == 94)
||(x_pointer == 98 && y_pointer == 94)
||(x_pointer == 99 && y_pointer == 94)
||(x_pointer == 100 && y_pointer == 94)
||(x_pointer == 101 && y_pointer == 94)
||(x_pointer == 102 && y_pointer == 94)
||(x_pointer == 103 && y_pointer == 94)
||(x_pointer == 104 && y_pointer == 94)
||(x_pointer == 105 && y_pointer == 94)
||(x_pointer == 106 && y_pointer == 94)
||(x_pointer == 107 && y_pointer == 94)
||(x_pointer == 108 && y_pointer == 94)
||(x_pointer == 109 && y_pointer == 94)
||(x_pointer == 110 && y_pointer == 94)
||(x_pointer == 111 && y_pointer == 94)
||(x_pointer == 112 && y_pointer == 94)
||(x_pointer == 113 && y_pointer == 94)
||(x_pointer == 114 && y_pointer == 94)
||(x_pointer == 115 && y_pointer == 94)
||(x_pointer == 116 && y_pointer == 94)
||(x_pointer == 117 && y_pointer == 94)
||(x_pointer == 118 && y_pointer == 94)
||(x_pointer == 119 && y_pointer == 94)
||(x_pointer == 120 && y_pointer == 94)
||(x_pointer == 36 && y_pointer == 95)
||(x_pointer == 37 && y_pointer == 95)
||(x_pointer == 38 && y_pointer == 95)
||(x_pointer == 39 && y_pointer == 95)
||(x_pointer == 40 && y_pointer == 95)
||(x_pointer == 41 && y_pointer == 95)
||(x_pointer == 42 && y_pointer == 95)
||(x_pointer == 43 && y_pointer == 95)
||(x_pointer == 44 && y_pointer == 95)
||(x_pointer == 45 && y_pointer == 95)
||(x_pointer == 46 && y_pointer == 95)
||(x_pointer == 47 && y_pointer == 95)
||(x_pointer == 48 && y_pointer == 95)
||(x_pointer == 49 && y_pointer == 95)
||(x_pointer == 50 && y_pointer == 95)
||(x_pointer == 51 && y_pointer == 95)
||(x_pointer == 52 && y_pointer == 95)
||(x_pointer == 53 && y_pointer == 95)
||(x_pointer == 54 && y_pointer == 95)
||(x_pointer == 55 && y_pointer == 95)
||(x_pointer == 56 && y_pointer == 95)
||(x_pointer == 57 && y_pointer == 95)
||(x_pointer == 58 && y_pointer == 95)
||(x_pointer == 59 && y_pointer == 95)
||(x_pointer == 60 && y_pointer == 95)
||(x_pointer == 67 && y_pointer == 95)
||(x_pointer == 68 && y_pointer == 95)
||(x_pointer == 69 && y_pointer == 95)
||(x_pointer == 70 && y_pointer == 95)
||(x_pointer == 71 && y_pointer == 95)
||(x_pointer == 72 && y_pointer == 95)
||(x_pointer == 73 && y_pointer == 95)
||(x_pointer == 74 && y_pointer == 95)
||(x_pointer == 75 && y_pointer == 95)
||(x_pointer == 76 && y_pointer == 95)
||(x_pointer == 77 && y_pointer == 95)
||(x_pointer == 78 && y_pointer == 95)
||(x_pointer == 79 && y_pointer == 95)
||(x_pointer == 80 && y_pointer == 95)
||(x_pointer == 81 && y_pointer == 95)
||(x_pointer == 82 && y_pointer == 95)
||(x_pointer == 83 && y_pointer == 95)
||(x_pointer == 84 && y_pointer == 95)
||(x_pointer == 85 && y_pointer == 95)
||(x_pointer == 86 && y_pointer == 95)
||(x_pointer == 87 && y_pointer == 95)
||(x_pointer == 88 && y_pointer == 95)
||(x_pointer == 89 && y_pointer == 95)
||(x_pointer == 96 && y_pointer == 95)
||(x_pointer == 97 && y_pointer == 95)
||(x_pointer == 98 && y_pointer == 95)
||(x_pointer == 99 && y_pointer == 95)
||(x_pointer == 100 && y_pointer == 95)
||(x_pointer == 101 && y_pointer == 95)
||(x_pointer == 102 && y_pointer == 95)
||(x_pointer == 103 && y_pointer == 95)
||(x_pointer == 104 && y_pointer == 95)
||(x_pointer == 105 && y_pointer == 95)
||(x_pointer == 106 && y_pointer == 95)
||(x_pointer == 107 && y_pointer == 95)
||(x_pointer == 108 && y_pointer == 95)
||(x_pointer == 109 && y_pointer == 95)
||(x_pointer == 110 && y_pointer == 95)
||(x_pointer == 111 && y_pointer == 95)
||(x_pointer == 112 && y_pointer == 95)
||(x_pointer == 113 && y_pointer == 95)
||(x_pointer == 114 && y_pointer == 95)
||(x_pointer == 115 && y_pointer == 95)
||(x_pointer == 116 && y_pointer == 95)
||(x_pointer == 117 && y_pointer == 95)
||(x_pointer == 118 && y_pointer == 95)
||(x_pointer == 119 && y_pointer == 95)
||(x_pointer == 120 && y_pointer == 95)
||(x_pointer == 36 && y_pointer == 96)
||(x_pointer == 37 && y_pointer == 96)
||(x_pointer == 38 && y_pointer == 96)
||(x_pointer == 39 && y_pointer == 96)
||(x_pointer == 40 && y_pointer == 96)
||(x_pointer == 41 && y_pointer == 96)
||(x_pointer == 42 && y_pointer == 96)
||(x_pointer == 43 && y_pointer == 96)
||(x_pointer == 44 && y_pointer == 96)
||(x_pointer == 45 && y_pointer == 96)
||(x_pointer == 46 && y_pointer == 96)
||(x_pointer == 47 && y_pointer == 96)
||(x_pointer == 48 && y_pointer == 96)
||(x_pointer == 49 && y_pointer == 96)
||(x_pointer == 50 && y_pointer == 96)
||(x_pointer == 51 && y_pointer == 96)
||(x_pointer == 52 && y_pointer == 96)
||(x_pointer == 53 && y_pointer == 96)
||(x_pointer == 54 && y_pointer == 96)
||(x_pointer == 55 && y_pointer == 96)
||(x_pointer == 56 && y_pointer == 96)
||(x_pointer == 57 && y_pointer == 96)
||(x_pointer == 58 && y_pointer == 96)
||(x_pointer == 59 && y_pointer == 96)
||(x_pointer == 60 && y_pointer == 96)
||(x_pointer == 67 && y_pointer == 96)
||(x_pointer == 68 && y_pointer == 96)
||(x_pointer == 69 && y_pointer == 96)
||(x_pointer == 70 && y_pointer == 96)
||(x_pointer == 71 && y_pointer == 96)
||(x_pointer == 72 && y_pointer == 96)
||(x_pointer == 73 && y_pointer == 96)
||(x_pointer == 74 && y_pointer == 96)
||(x_pointer == 75 && y_pointer == 96)
||(x_pointer == 76 && y_pointer == 96)
||(x_pointer == 77 && y_pointer == 96)
||(x_pointer == 78 && y_pointer == 96)
||(x_pointer == 79 && y_pointer == 96)
||(x_pointer == 80 && y_pointer == 96)
||(x_pointer == 81 && y_pointer == 96)
||(x_pointer == 82 && y_pointer == 96)
||(x_pointer == 83 && y_pointer == 96)
||(x_pointer == 84 && y_pointer == 96)
||(x_pointer == 85 && y_pointer == 96)
||(x_pointer == 86 && y_pointer == 96)
||(x_pointer == 87 && y_pointer == 96)
||(x_pointer == 88 && y_pointer == 96)
||(x_pointer == 89 && y_pointer == 96)
||(x_pointer == 96 && y_pointer == 96)
||(x_pointer == 97 && y_pointer == 96)
||(x_pointer == 98 && y_pointer == 96)
||(x_pointer == 99 && y_pointer == 96)
||(x_pointer == 100 && y_pointer == 96)
||(x_pointer == 101 && y_pointer == 96)
||(x_pointer == 102 && y_pointer == 96)
||(x_pointer == 103 && y_pointer == 96)
||(x_pointer == 104 && y_pointer == 96)
||(x_pointer == 105 && y_pointer == 96)
||(x_pointer == 106 && y_pointer == 96)
||(x_pointer == 107 && y_pointer == 96)
||(x_pointer == 108 && y_pointer == 96)
||(x_pointer == 109 && y_pointer == 96)
||(x_pointer == 110 && y_pointer == 96)
||(x_pointer == 111 && y_pointer == 96)
||(x_pointer == 112 && y_pointer == 96)
||(x_pointer == 113 && y_pointer == 96)
||(x_pointer == 114 && y_pointer == 96)
||(x_pointer == 115 && y_pointer == 96)
||(x_pointer == 116 && y_pointer == 96)
||(x_pointer == 117 && y_pointer == 96)
||(x_pointer == 118 && y_pointer == 96)
||(x_pointer == 119 && y_pointer == 96)
||(x_pointer == 120 && y_pointer == 96)
||(x_pointer == 36 && y_pointer == 97)
||(x_pointer == 37 && y_pointer == 97)
||(x_pointer == 38 && y_pointer == 97)
||(x_pointer == 39 && y_pointer == 97)
||(x_pointer == 40 && y_pointer == 97)
||(x_pointer == 41 && y_pointer == 97)
||(x_pointer == 42 && y_pointer == 97)
||(x_pointer == 43 && y_pointer == 97)
||(x_pointer == 44 && y_pointer == 97)
||(x_pointer == 45 && y_pointer == 97)
||(x_pointer == 46 && y_pointer == 97)
||(x_pointer == 47 && y_pointer == 97)
||(x_pointer == 48 && y_pointer == 97)
||(x_pointer == 49 && y_pointer == 97)
||(x_pointer == 50 && y_pointer == 97)
||(x_pointer == 51 && y_pointer == 97)
||(x_pointer == 52 && y_pointer == 97)
||(x_pointer == 53 && y_pointer == 97)
||(x_pointer == 54 && y_pointer == 97)
||(x_pointer == 55 && y_pointer == 97)
||(x_pointer == 56 && y_pointer == 97)
||(x_pointer == 57 && y_pointer == 97)
||(x_pointer == 58 && y_pointer == 97)
||(x_pointer == 59 && y_pointer == 97)
||(x_pointer == 60 && y_pointer == 97)
||(x_pointer == 67 && y_pointer == 97)
||(x_pointer == 68 && y_pointer == 97)
||(x_pointer == 69 && y_pointer == 97)
||(x_pointer == 70 && y_pointer == 97)
||(x_pointer == 71 && y_pointer == 97)
||(x_pointer == 72 && y_pointer == 97)
||(x_pointer == 73 && y_pointer == 97)
||(x_pointer == 74 && y_pointer == 97)
||(x_pointer == 75 && y_pointer == 97)
||(x_pointer == 76 && y_pointer == 97)
||(x_pointer == 77 && y_pointer == 97)
||(x_pointer == 78 && y_pointer == 97)
||(x_pointer == 79 && y_pointer == 97)
||(x_pointer == 80 && y_pointer == 97)
||(x_pointer == 81 && y_pointer == 97)
||(x_pointer == 82 && y_pointer == 97)
||(x_pointer == 83 && y_pointer == 97)
||(x_pointer == 84 && y_pointer == 97)
||(x_pointer == 85 && y_pointer == 97)
||(x_pointer == 86 && y_pointer == 97)
||(x_pointer == 87 && y_pointer == 97)
||(x_pointer == 88 && y_pointer == 97)
||(x_pointer == 89 && y_pointer == 97)
||(x_pointer == 96 && y_pointer == 97)
||(x_pointer == 97 && y_pointer == 97)
||(x_pointer == 98 && y_pointer == 97)
||(x_pointer == 99 && y_pointer == 97)
||(x_pointer == 100 && y_pointer == 97)
||(x_pointer == 101 && y_pointer == 97)
||(x_pointer == 102 && y_pointer == 97)
||(x_pointer == 103 && y_pointer == 97)
||(x_pointer == 104 && y_pointer == 97)
||(x_pointer == 105 && y_pointer == 97)
||(x_pointer == 106 && y_pointer == 97)
||(x_pointer == 107 && y_pointer == 97)
||(x_pointer == 108 && y_pointer == 97)
||(x_pointer == 109 && y_pointer == 97)
||(x_pointer == 110 && y_pointer == 97)
||(x_pointer == 111 && y_pointer == 97)
||(x_pointer == 112 && y_pointer == 97)
||(x_pointer == 113 && y_pointer == 97)
||(x_pointer == 114 && y_pointer == 97)
||(x_pointer == 115 && y_pointer == 97)
||(x_pointer == 116 && y_pointer == 97)
||(x_pointer == 117 && y_pointer == 97)
||(x_pointer == 118 && y_pointer == 97)
||(x_pointer == 119 && y_pointer == 97)
||(x_pointer == 120 && y_pointer == 97));
endmodule