module game_text_setter(clk, score, ingame, main_difficulty, x_pointer, y_pointer, game_text);
   input ingame;
	input [3:0] main_difficulty;
   input clk;
   input [7:0]x_pointer;
	input [6:0]y_pointer;
	input [12:0] score;
	output reg game_text; // check if the pixel is the menu's text.
	

	
	reg [3:0] units_digit_score;
	reg [3:0] tens_digit_score;
	reg [3:0] hundreds_digit_score;
	
	
	always@(posedge clk)begin
		units_digit_score <= score % 10;
	   tens_digit_score <= ((score - (score % 10)) / 10) % 10;
		hundreds_digit_score <= (score - (score % 10) - 	(10 * ((score - (score % 10)) / 10) % 10)) / 100;
	end
	

	//menu's normal text
	always@(posedge clk)
	begin
		if (ingame)
			 begin
			 if (main_texts
			     ||easy
				  ||normal
				  ||hard
				  ||units_digit_0
				  ||units_digit_1
				  ||units_digit_2
				  ||units_digit_3
				  ||units_digit_4
				  ||units_digit_5
				  ||units_digit_6
				  ||units_digit_7
				  ||units_digit_8
				  ||units_digit_9
				  )
				 game_text <= 1'b1;
			 else
				 game_text <= 1'b0;
			 end
	end
	
	
	
	
	// wires for main texts
	wire main_texts = 
	(x_pointer == 5 && y_pointer == 114)
||(x_pointer == 6 && y_pointer == 114)
||(x_pointer == 7 && y_pointer == 114)
||(x_pointer == 8 && y_pointer == 114)
||(x_pointer == 10 && y_pointer == 114)
||(x_pointer == 11 && y_pointer == 114)
||(x_pointer == 12 && y_pointer == 114)
||(x_pointer == 13 && y_pointer == 114)
||(x_pointer == 15 && y_pointer == 114)
||(x_pointer == 16 && y_pointer == 114)
||(x_pointer == 17 && y_pointer == 114)
||(x_pointer == 18 && y_pointer == 114)
||(x_pointer == 20 && y_pointer == 114)
||(x_pointer == 21 && y_pointer == 114)
||(x_pointer == 22 && y_pointer == 114)
||(x_pointer == 23 && y_pointer == 114)
||(x_pointer == 25 && y_pointer == 114)
||(x_pointer == 26 && y_pointer == 114)
||(x_pointer == 27 && y_pointer == 114)
||(x_pointer == 28 && y_pointer == 114)
||(x_pointer == 48 && y_pointer == 114)
||(x_pointer == 51 && y_pointer == 114)
||(x_pointer == 53 && y_pointer == 114)
||(x_pointer == 55 && y_pointer == 114)
||(x_pointer == 56 && y_pointer == 114)
||(x_pointer == 57 && y_pointer == 114)
||(x_pointer == 58 && y_pointer == 114)
||(x_pointer == 60 && y_pointer == 114)
||(x_pointer == 61 && y_pointer == 114)
||(x_pointer == 62 && y_pointer == 114)
||(x_pointer == 63 && y_pointer == 114)
||(x_pointer == 65 && y_pointer == 114)
||(x_pointer == 66 && y_pointer == 114)
||(x_pointer == 67 && y_pointer == 114)
||(x_pointer == 68 && y_pointer == 114)
||(x_pointer == 70 && y_pointer == 114)
||(x_pointer == 71 && y_pointer == 114)
||(x_pointer == 72 && y_pointer == 114)
||(x_pointer == 73 && y_pointer == 114)
||(x_pointer == 75 && y_pointer == 114)
||(x_pointer == 76 && y_pointer == 114)
||(x_pointer == 77 && y_pointer == 114)
||(x_pointer == 78 && y_pointer == 114)
||(x_pointer == 99 && y_pointer == 114)
||(x_pointer == 103 && y_pointer == 114)
||(x_pointer == 104 && y_pointer == 114)
||(x_pointer == 105 && y_pointer == 114)
||(x_pointer == 106 && y_pointer == 114)
||(x_pointer == 108 && y_pointer == 114)
||(x_pointer == 110 && y_pointer == 114)
||(x_pointer == 112 && y_pointer == 114)
||(x_pointer == 113 && y_pointer == 114)
||(x_pointer == 114 && y_pointer == 114)
||(x_pointer == 115 && y_pointer == 114)
||(x_pointer == 117 && y_pointer == 114)
||(x_pointer == 5 && y_pointer == 115)
||(x_pointer == 10 && y_pointer == 115)
||(x_pointer == 15 && y_pointer == 115)
||(x_pointer == 18 && y_pointer == 115)
||(x_pointer == 20 && y_pointer == 115)
||(x_pointer == 23 && y_pointer == 115)
||(x_pointer == 25 && y_pointer == 115)
||(x_pointer == 48 && y_pointer == 115)
||(x_pointer == 51 && y_pointer == 115)
||(x_pointer == 53 && y_pointer == 115)
||(x_pointer == 55 && y_pointer == 115)
||(x_pointer == 60 && y_pointer == 115)
||(x_pointer == 65 && y_pointer == 115)
||(x_pointer == 68 && y_pointer == 115)
||(x_pointer == 70 && y_pointer == 115)
||(x_pointer == 73 && y_pointer == 115)
||(x_pointer == 75 && y_pointer == 115)
||(x_pointer == 99 && y_pointer == 115)
||(x_pointer == 103 && y_pointer == 115)
||(x_pointer == 108 && y_pointer == 115)
||(x_pointer == 110 && y_pointer == 115)
||(x_pointer == 112 && y_pointer == 115)
||(x_pointer == 117 && y_pointer == 115)
||(x_pointer == 5 && y_pointer == 116)
||(x_pointer == 6 && y_pointer == 116)
||(x_pointer == 7 && y_pointer == 116)
||(x_pointer == 8 && y_pointer == 116)
||(x_pointer == 10 && y_pointer == 116)
||(x_pointer == 15 && y_pointer == 116)
||(x_pointer == 18 && y_pointer == 116)
||(x_pointer == 20 && y_pointer == 116)
||(x_pointer == 21 && y_pointer == 116)
||(x_pointer == 22 && y_pointer == 116)
||(x_pointer == 23 && y_pointer == 116)
||(x_pointer == 25 && y_pointer == 116)
||(x_pointer == 26 && y_pointer == 116)
||(x_pointer == 27 && y_pointer == 116)
||(x_pointer == 28 && y_pointer == 116)
||(x_pointer == 48 && y_pointer == 116)
||(x_pointer == 49 && y_pointer == 116)
||(x_pointer == 50 && y_pointer == 116)
||(x_pointer == 51 && y_pointer == 116)
||(x_pointer == 53 && y_pointer == 116)
||(x_pointer == 55 && y_pointer == 116)
||(x_pointer == 56 && y_pointer == 116)
||(x_pointer == 57 && y_pointer == 116)
||(x_pointer == 58 && y_pointer == 116)
||(x_pointer == 60 && y_pointer == 116)
||(x_pointer == 65 && y_pointer == 116)
||(x_pointer == 68 && y_pointer == 116)
||(x_pointer == 70 && y_pointer == 116)
||(x_pointer == 71 && y_pointer == 116)
||(x_pointer == 72 && y_pointer == 116)
||(x_pointer == 73 && y_pointer == 116)
||(x_pointer == 75 && y_pointer == 116)
||(x_pointer == 76 && y_pointer == 116)
||(x_pointer == 77 && y_pointer == 116)
||(x_pointer == 78 && y_pointer == 116)
||(x_pointer == 99 && y_pointer == 116)
||(x_pointer == 103 && y_pointer == 116)
||(x_pointer == 104 && y_pointer == 116)
||(x_pointer == 105 && y_pointer == 116)
||(x_pointer == 106 && y_pointer == 116)
||(x_pointer == 108 && y_pointer == 116)
||(x_pointer == 110 && y_pointer == 116)
||(x_pointer == 112 && y_pointer == 116)
||(x_pointer == 113 && y_pointer == 116)
||(x_pointer == 114 && y_pointer == 116)
||(x_pointer == 115 && y_pointer == 116)
||(x_pointer == 117 && y_pointer == 116)
||(x_pointer == 8 && y_pointer == 117)
||(x_pointer == 10 && y_pointer == 117)
||(x_pointer == 15 && y_pointer == 117)
||(x_pointer == 18 && y_pointer == 117)
||(x_pointer == 20 && y_pointer == 117)
||(x_pointer == 21 && y_pointer == 117)
||(x_pointer == 25 && y_pointer == 117)
||(x_pointer == 48 && y_pointer == 117)
||(x_pointer == 51 && y_pointer == 117)
||(x_pointer == 53 && y_pointer == 117)
||(x_pointer == 58 && y_pointer == 117)
||(x_pointer == 60 && y_pointer == 117)
||(x_pointer == 65 && y_pointer == 117)
||(x_pointer == 68 && y_pointer == 117)
||(x_pointer == 70 && y_pointer == 117)
||(x_pointer == 71 && y_pointer == 117)
||(x_pointer == 75 && y_pointer == 117)
||(x_pointer == 99 && y_pointer == 117)
||(x_pointer == 103 && y_pointer == 117)
||(x_pointer == 108 && y_pointer == 117)
||(x_pointer == 110 && y_pointer == 117)
||(x_pointer == 112 && y_pointer == 117)
||(x_pointer == 117 && y_pointer == 117)
||(x_pointer == 5 && y_pointer == 118)
||(x_pointer == 6 && y_pointer == 118)
||(x_pointer == 7 && y_pointer == 118)
||(x_pointer == 8 && y_pointer == 118)
||(x_pointer == 10 && y_pointer == 118)
||(x_pointer == 11 && y_pointer == 118)
||(x_pointer == 12 && y_pointer == 118)
||(x_pointer == 13 && y_pointer == 118)
||(x_pointer == 15 && y_pointer == 118)
||(x_pointer == 16 && y_pointer == 118)
||(x_pointer == 17 && y_pointer == 118)
||(x_pointer == 18 && y_pointer == 118)
||(x_pointer == 20 && y_pointer == 118)
||(x_pointer == 22 && y_pointer == 118)
||(x_pointer == 23 && y_pointer == 118)
||(x_pointer == 25 && y_pointer == 118)
||(x_pointer == 26 && y_pointer == 118)
||(x_pointer == 27 && y_pointer == 118)
||(x_pointer == 28 && y_pointer == 118)
||(x_pointer == 48 && y_pointer == 118)
||(x_pointer == 51 && y_pointer == 118)
||(x_pointer == 53 && y_pointer == 118)
||(x_pointer == 55 && y_pointer == 118)
||(x_pointer == 56 && y_pointer == 118)
||(x_pointer == 57 && y_pointer == 118)
||(x_pointer == 58 && y_pointer == 118)
||(x_pointer == 60 && y_pointer == 118)
||(x_pointer == 61 && y_pointer == 118)
||(x_pointer == 62 && y_pointer == 118)
||(x_pointer == 63 && y_pointer == 118)
||(x_pointer == 65 && y_pointer == 118)
||(x_pointer == 66 && y_pointer == 118)
||(x_pointer == 67 && y_pointer == 118)
||(x_pointer == 68 && y_pointer == 118)
||(x_pointer == 70 && y_pointer == 118)
||(x_pointer == 72 && y_pointer == 118)
||(x_pointer == 73 && y_pointer == 118)
||(x_pointer == 75 && y_pointer == 118)
||(x_pointer == 76 && y_pointer == 118)
||(x_pointer == 77 && y_pointer == 118)
||(x_pointer == 78 && y_pointer == 118)
||(x_pointer == 99 && y_pointer == 118)
||(x_pointer == 100 && y_pointer == 118)
||(x_pointer == 101 && y_pointer == 118)
||(x_pointer == 103 && y_pointer == 118)
||(x_pointer == 104 && y_pointer == 118)
||(x_pointer == 105 && y_pointer == 118)
||(x_pointer == 106 && y_pointer == 118)
||(x_pointer == 109 && y_pointer == 118)
||(x_pointer == 112 && y_pointer == 118)
||(x_pointer == 113 && y_pointer == 118)
||(x_pointer == 114 && y_pointer == 118)
||(x_pointer == 115 && y_pointer == 118)
||(x_pointer == 117 && y_pointer == 118)
||(x_pointer == 118 && y_pointer == 118)
||(x_pointer == 119 && y_pointer == 118);

   wire easy = 
	main_difficulty == 4'd1 && ((x_pointer == 134 && y_pointer == 114)
||(x_pointer == 137 && y_pointer == 114)
||(x_pointer == 140 && y_pointer == 114)
||(x_pointer == 141 && y_pointer == 114)
||(x_pointer == 144 && y_pointer == 114)
||(x_pointer == 145 && y_pointer == 114)
||(x_pointer == 146 && y_pointer == 114)
||(x_pointer == 147 && y_pointer == 114)
||(x_pointer == 149 && y_pointer == 114)
||(x_pointer == 150 && y_pointer == 114)
||(x_pointer == 151 && y_pointer == 114)
||(x_pointer == 134 && y_pointer == 115)
||(x_pointer == 137 && y_pointer == 115)
||(x_pointer == 139 && y_pointer == 115)
||(x_pointer == 142 && y_pointer == 115)
||(x_pointer == 144 && y_pointer == 115)
||(x_pointer == 147 && y_pointer == 115)
||(x_pointer == 149 && y_pointer == 115)
||(x_pointer == 152 && y_pointer == 115)
||(x_pointer == 134 && y_pointer == 116)
||(x_pointer == 135 && y_pointer == 116)
||(x_pointer == 136 && y_pointer == 116)
||(x_pointer == 137 && y_pointer == 116)
||(x_pointer == 139 && y_pointer == 116)
||(x_pointer == 140 && y_pointer == 116)
||(x_pointer == 141 && y_pointer == 116)
||(x_pointer == 142 && y_pointer == 116)
||(x_pointer == 144 && y_pointer == 116)
||(x_pointer == 145 && y_pointer == 116)
||(x_pointer == 146 && y_pointer == 116)
||(x_pointer == 147 && y_pointer == 116)
||(x_pointer == 149 && y_pointer == 116)
||(x_pointer == 152 && y_pointer == 116)
||(x_pointer == 134 && y_pointer == 117)
||(x_pointer == 137 && y_pointer == 117)
||(x_pointer == 139 && y_pointer == 117)
||(x_pointer == 142 && y_pointer == 117)
||(x_pointer == 144 && y_pointer == 117)
||(x_pointer == 145 && y_pointer == 117)
||(x_pointer == 149 && y_pointer == 117)
||(x_pointer == 152 && y_pointer == 117)
||(x_pointer == 134 && y_pointer == 118)
||(x_pointer == 137 && y_pointer == 118)
||(x_pointer == 139 && y_pointer == 118)
||(x_pointer == 142 && y_pointer == 118)
||(x_pointer == 144 && y_pointer == 118)
||(x_pointer == 146 && y_pointer == 118)
||(x_pointer == 147 && y_pointer == 118)
||(x_pointer == 149 && y_pointer == 118)
||(x_pointer == 150 && y_pointer == 118)
||(x_pointer == 151 && y_pointer == 118));
	
	wire normal = 
	main_difficulty == 4'd2 && ((x_pointer == 128 && y_pointer == 114)
||(x_pointer == 132 && y_pointer == 114)
||(x_pointer == 134 && y_pointer == 114)
||(x_pointer == 135 && y_pointer == 114)
||(x_pointer == 136 && y_pointer == 114)
||(x_pointer == 137 && y_pointer == 114)
||(x_pointer == 139 && y_pointer == 114)
||(x_pointer == 140 && y_pointer == 114)
||(x_pointer == 141 && y_pointer == 114)
||(x_pointer == 142 && y_pointer == 114)
||(x_pointer == 144 && y_pointer == 114)
||(x_pointer == 148 && y_pointer == 114)
||(x_pointer == 151 && y_pointer == 114)
||(x_pointer == 152 && y_pointer == 114)
||(x_pointer == 155 && y_pointer == 114)
||(x_pointer == 128 && y_pointer == 115)
||(x_pointer == 129 && y_pointer == 115)
||(x_pointer == 132 && y_pointer == 115)
||(x_pointer == 134 && y_pointer == 115)
||(x_pointer == 137 && y_pointer == 115)
||(x_pointer == 139 && y_pointer == 115)
||(x_pointer == 142 && y_pointer == 115)
||(x_pointer == 144 && y_pointer == 115)
||(x_pointer == 145 && y_pointer == 115)
||(x_pointer == 147 && y_pointer == 115)
||(x_pointer == 148 && y_pointer == 115)
||(x_pointer == 150 && y_pointer == 115)
||(x_pointer == 153 && y_pointer == 115)
||(x_pointer == 155 && y_pointer == 115)
||(x_pointer == 128 && y_pointer == 116)
||(x_pointer == 130 && y_pointer == 116)
||(x_pointer == 132 && y_pointer == 116)
||(x_pointer == 134 && y_pointer == 116)
||(x_pointer == 137 && y_pointer == 116)
||(x_pointer == 139 && y_pointer == 116)
||(x_pointer == 140 && y_pointer == 116)
||(x_pointer == 141 && y_pointer == 116)
||(x_pointer == 142 && y_pointer == 116)
||(x_pointer == 144 && y_pointer == 116)
||(x_pointer == 146 && y_pointer == 116)
||(x_pointer == 148 && y_pointer == 116)
||(x_pointer == 150 && y_pointer == 116)
||(x_pointer == 151 && y_pointer == 116)
||(x_pointer == 152 && y_pointer == 116)
||(x_pointer == 153 && y_pointer == 116)
||(x_pointer == 155 && y_pointer == 116)
||(x_pointer == 128 && y_pointer == 117)
||(x_pointer == 131 && y_pointer == 117)
||(x_pointer == 132 && y_pointer == 117)
||(x_pointer == 134 && y_pointer == 117)
||(x_pointer == 137 && y_pointer == 117)
||(x_pointer == 139 && y_pointer == 117)
||(x_pointer == 140 && y_pointer == 117)
||(x_pointer == 144 && y_pointer == 117)
||(x_pointer == 146 && y_pointer == 117)
||(x_pointer == 148 && y_pointer == 117)
||(x_pointer == 150 && y_pointer == 117)
||(x_pointer == 153 && y_pointer == 117)
||(x_pointer == 155 && y_pointer == 117)
||(x_pointer == 128 && y_pointer == 118)
||(x_pointer == 132 && y_pointer == 118)
||(x_pointer == 134 && y_pointer == 118)
||(x_pointer == 135 && y_pointer == 118)
||(x_pointer == 136 && y_pointer == 118)
||(x_pointer == 137 && y_pointer == 118)
||(x_pointer == 139 && y_pointer == 118)
||(x_pointer == 141 && y_pointer == 118)
||(x_pointer == 142 && y_pointer == 118)
||(x_pointer == 144 && y_pointer == 118)
||(x_pointer == 148 && y_pointer == 118)
||(x_pointer == 150 && y_pointer == 118)
||(x_pointer == 153 && y_pointer == 118)
||(x_pointer == 155 && y_pointer == 118)
||(x_pointer == 156 && y_pointer == 118)
||(x_pointer == 157 && y_pointer == 118));
	
	wire hard = 
	main_difficulty == 4'd4 && ((x_pointer == 134 && y_pointer == 114)
||(x_pointer == 135 && y_pointer == 114)
||(x_pointer == 136 && y_pointer == 114)
||(x_pointer == 137 && y_pointer == 114)
||(x_pointer == 140 && y_pointer == 114)
||(x_pointer == 141 && y_pointer == 114)
||(x_pointer == 144 && y_pointer == 114)
||(x_pointer == 145 && y_pointer == 114)
||(x_pointer == 146 && y_pointer == 114)
||(x_pointer == 147 && y_pointer == 114)
||(x_pointer == 149 && y_pointer == 114)
||(x_pointer == 151 && y_pointer == 114)
||(x_pointer == 134 && y_pointer == 115)
||(x_pointer == 139 && y_pointer == 115)
||(x_pointer == 142 && y_pointer == 115)
||(x_pointer == 144 && y_pointer == 115)
||(x_pointer == 149 && y_pointer == 115)
||(x_pointer == 151 && y_pointer == 115)
||(x_pointer == 134 && y_pointer == 116)
||(x_pointer == 135 && y_pointer == 116)
||(x_pointer == 136 && y_pointer == 116)
||(x_pointer == 137 && y_pointer == 116)
||(x_pointer == 139 && y_pointer == 116)
||(x_pointer == 140 && y_pointer == 116)
||(x_pointer == 141 && y_pointer == 116)
||(x_pointer == 142 && y_pointer == 116)
||(x_pointer == 144 && y_pointer == 116)
||(x_pointer == 145 && y_pointer == 116)
||(x_pointer == 146 && y_pointer == 116)
||(x_pointer == 147 && y_pointer == 116)
||(x_pointer == 149 && y_pointer == 116)
||(x_pointer == 151 && y_pointer == 116)
||(x_pointer == 134 && y_pointer == 117)
||(x_pointer == 139 && y_pointer == 117)
||(x_pointer == 142 && y_pointer == 117)
||(x_pointer == 147 && y_pointer == 117)
||(x_pointer == 150 && y_pointer == 117)
||(x_pointer == 134 && y_pointer == 118)
||(x_pointer == 135 && y_pointer == 118)
||(x_pointer == 136 && y_pointer == 118)
||(x_pointer == 137 && y_pointer == 118)
||(x_pointer == 139 && y_pointer == 118)
||(x_pointer == 142 && y_pointer == 118)
||(x_pointer == 144 && y_pointer == 118)
||(x_pointer == 145 && y_pointer == 118)
||(x_pointer == 146 && y_pointer == 118)
||(x_pointer == 147 && y_pointer == 118)
||(x_pointer == 150 && y_pointer == 118));
   wire units_digit_0 = units_digit_score == 0 && ((x_pointer == 42 && y_pointer == 114)
||(x_pointer == 43 && y_pointer == 114)
||(x_pointer == 44 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 114)
||(x_pointer == 42 && y_pointer == 115)
||(x_pointer == 45 && y_pointer == 115)
||(x_pointer == 42 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 116)
||(x_pointer == 42 && y_pointer == 117)
||(x_pointer == 45 && y_pointer == 117)
||(x_pointer == 42 && y_pointer == 118)
||(x_pointer == 43 && y_pointer == 118)
||(x_pointer == 44 && y_pointer == 118)
||(x_pointer == 45 && y_pointer == 118));
	wire units_digit_1 = units_digit_score == 1 && ((x_pointer == 45 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 115)
||(x_pointer == 45 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 117)
||(x_pointer == 45 && y_pointer == 118));
   wire units_digit_2 = units_digit_score == 2 && ((x_pointer == 42 && y_pointer == 114)
||(x_pointer == 43 && y_pointer == 114)
||(x_pointer == 44 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 115)
||(x_pointer == 42 && y_pointer == 116)
||(x_pointer == 43 && y_pointer == 116)
||(x_pointer == 44 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 116)
||(x_pointer == 42 && y_pointer == 117)
||(x_pointer == 42 && y_pointer == 118)
||(x_pointer == 43 && y_pointer == 118)
||(x_pointer == 44 && y_pointer == 118)
||(x_pointer == 45 && y_pointer == 118));
	wire units_digit_3 = units_digit_score == 3 && ((x_pointer == 42 && y_pointer == 114)
||(x_pointer == 43 && y_pointer == 114)
||(x_pointer == 44 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 115)
||(x_pointer == 42 && y_pointer == 116)
||(x_pointer == 43 && y_pointer == 116)
||(x_pointer == 44 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 117)
||(x_pointer == 42 && y_pointer == 118)
||(x_pointer == 43 && y_pointer == 118)
||(x_pointer == 44 && y_pointer == 118)
||(x_pointer == 45 && y_pointer == 118));
	wire units_digit_4 = units_digit_score == 4 && ((x_pointer == 42 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 114)
||(x_pointer == 42 && y_pointer == 115)
||(x_pointer == 45 && y_pointer == 115)
||(x_pointer == 42 && y_pointer == 116)
||(x_pointer == 43 && y_pointer == 116)
||(x_pointer == 44 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 117)
||(x_pointer == 45 && y_pointer == 118));
	wire units_digit_5 = units_digit_score == 5 && ((x_pointer == 42 && y_pointer == 114)
||(x_pointer == 43 && y_pointer == 114)
||(x_pointer == 44 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 114)
||(x_pointer == 42 && y_pointer == 115)
||(x_pointer == 42 && y_pointer == 116)
||(x_pointer == 43 && y_pointer == 116)
||(x_pointer == 44 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 117)
||(x_pointer == 42 && y_pointer == 118)
||(x_pointer == 43 && y_pointer == 118)
||(x_pointer == 44 && y_pointer == 118)
||(x_pointer == 45 && y_pointer == 118));
	wire units_digit_6 = units_digit_score == 6 && ((x_pointer == 42 && y_pointer == 114)
||(x_pointer == 43 && y_pointer == 114)
||(x_pointer == 44 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 114)
||(x_pointer == 42 && y_pointer == 115)
||(x_pointer == 42 && y_pointer == 116)
||(x_pointer == 43 && y_pointer == 116)
||(x_pointer == 44 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 116)
||(x_pointer == 42 && y_pointer == 117)
||(x_pointer == 45 && y_pointer == 117)
||(x_pointer == 42 && y_pointer == 118)
||(x_pointer == 43 && y_pointer == 118)
||(x_pointer == 44 && y_pointer == 118)
||(x_pointer == 45 && y_pointer == 118));
	wire units_digit_7 = units_digit_score == 7 && ((x_pointer == 42 && y_pointer == 114)
||(x_pointer == 43 && y_pointer == 114)
||(x_pointer == 44 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 115)
||(x_pointer == 45 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 117)
||(x_pointer == 45 && y_pointer == 118));
	wire units_digit_8 = units_digit_score == 8 && (
	(x_pointer == 42 && y_pointer == 114)
||(x_pointer == 43 && y_pointer == 114)
||(x_pointer == 44 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 114)
||(x_pointer == 42 && y_pointer == 115)
||(x_pointer == 45 && y_pointer == 115)
||(x_pointer == 42 && y_pointer == 116)
||(x_pointer == 43 && y_pointer == 116)
||(x_pointer == 44 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 116)
||(x_pointer == 42 && y_pointer == 117)
||(x_pointer == 45 && y_pointer == 117)
||(x_pointer == 42 && y_pointer == 118)
||(x_pointer == 43 && y_pointer == 118)
||(x_pointer == 44 && y_pointer == 118)
||(x_pointer == 45 && y_pointer == 118)
	);
	wire units_digit_9 = units_digit_score == 9 && ((x_pointer == 42 && y_pointer == 114)
||(x_pointer == 43 && y_pointer == 114)
||(x_pointer == 44 && y_pointer == 114)
||(x_pointer == 45 && y_pointer == 114)
||(x_pointer == 42 && y_pointer == 115)
||(x_pointer == 45 && y_pointer == 115)
||(x_pointer == 42 && y_pointer == 116)
||(x_pointer == 43 && y_pointer == 116)
||(x_pointer == 44 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 116)
||(x_pointer == 45 && y_pointer == 117)
||(x_pointer == 42 && y_pointer == 118)
||(x_pointer == 43 && y_pointer == 118)
||(x_pointer == 44 && y_pointer == 118)
||(x_pointer == 45 && y_pointer == 118));
endmodule