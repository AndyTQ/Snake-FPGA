module game_barrier_setter(clk, ingame, current_level, x_pointer, y_pointer, barrier);
   input ingame;
	input [3:0] current_level;
   input clk;
   input [7:0]x_pointer;
	input [6:0]y_pointer;
	output reg barrier; 

	always@(posedge clk)
	begin
		if (ingame)
			 begin
			 if (barrier_pixel_0 
			 || barrier_pixel_1 
			 || barrier_pixel_2
			 || barrier_pixel_3
			 || barrier_pixel_4
			 || barrier_pixel_5
			 || barrier_pixel_6
			 || barrier_pixel_7)
				 barrier <= 1'b1;
			 else
				 barrier <= 1'b0;
			 end
	end
	wire barrier_pixel_0 = 1'b0;
	wire barrier_pixel_1 = current_level == 1 && ((x_pointer == 29 && y_pointer == 53)
||(x_pointer == 30 && y_pointer == 53)
||(x_pointer == 31 && y_pointer == 53)
||(x_pointer == 32 && y_pointer == 53)
||(x_pointer == 33 && y_pointer == 53)
||(x_pointer == 34 && y_pointer == 53)
||(x_pointer == 35 && y_pointer == 53)
||(x_pointer == 36 && y_pointer == 53)
||(x_pointer == 37 && y_pointer == 53)
||(x_pointer == 38 && y_pointer == 53)
||(x_pointer == 39 && y_pointer == 53)
||(x_pointer == 40 && y_pointer == 53)
||(x_pointer == 41 && y_pointer == 53)
||(x_pointer == 42 && y_pointer == 53)
||(x_pointer == 43 && y_pointer == 53)
||(x_pointer == 44 && y_pointer == 53)
||(x_pointer == 45 && y_pointer == 53)
||(x_pointer == 46 && y_pointer == 53)
||(x_pointer == 47 && y_pointer == 53)
||(x_pointer == 48 && y_pointer == 53)
||(x_pointer == 49 && y_pointer == 53)
||(x_pointer == 50 && y_pointer == 53)
||(x_pointer == 51 && y_pointer == 53)
||(x_pointer == 52 && y_pointer == 53)
||(x_pointer == 53 && y_pointer == 53)
||(x_pointer == 54 && y_pointer == 53)
||(x_pointer == 55 && y_pointer == 53)
||(x_pointer == 56 && y_pointer == 53)
||(x_pointer == 57 && y_pointer == 53)
||(x_pointer == 58 && y_pointer == 53)
||(x_pointer == 59 && y_pointer == 53)
||(x_pointer == 60 && y_pointer == 53)
||(x_pointer == 61 && y_pointer == 53)
||(x_pointer == 62 && y_pointer == 53)
||(x_pointer == 63 && y_pointer == 53)
||(x_pointer == 64 && y_pointer == 53)
||(x_pointer == 65 && y_pointer == 53)
||(x_pointer == 66 && y_pointer == 53)
||(x_pointer == 67 && y_pointer == 53)
||(x_pointer == 92 && y_pointer == 53)
||(x_pointer == 93 && y_pointer == 53)
||(x_pointer == 94 && y_pointer == 53)
||(x_pointer == 95 && y_pointer == 53)
||(x_pointer == 96 && y_pointer == 53)
||(x_pointer == 97 && y_pointer == 53)
||(x_pointer == 98 && y_pointer == 53)
||(x_pointer == 99 && y_pointer == 53)
||(x_pointer == 100 && y_pointer == 53)
||(x_pointer == 101 && y_pointer == 53)
||(x_pointer == 102 && y_pointer == 53)
||(x_pointer == 103 && y_pointer == 53)
||(x_pointer == 104 && y_pointer == 53)
||(x_pointer == 105 && y_pointer == 53)
||(x_pointer == 106 && y_pointer == 53)
||(x_pointer == 107 && y_pointer == 53)
||(x_pointer == 108 && y_pointer == 53)
||(x_pointer == 109 && y_pointer == 53)
||(x_pointer == 110 && y_pointer == 53)
||(x_pointer == 111 && y_pointer == 53)
||(x_pointer == 112 && y_pointer == 53)
||(x_pointer == 113 && y_pointer == 53)
||(x_pointer == 114 && y_pointer == 53)
||(x_pointer == 115 && y_pointer == 53)
||(x_pointer == 116 && y_pointer == 53)
||(x_pointer == 117 && y_pointer == 53)
||(x_pointer == 118 && y_pointer == 53)
||(x_pointer == 119 && y_pointer == 53)
||(x_pointer == 120 && y_pointer == 53)
||(x_pointer == 121 && y_pointer == 53)
||(x_pointer == 122 && y_pointer == 53)
||(x_pointer == 123 && y_pointer == 53)
||(x_pointer == 124 && y_pointer == 53)
||(x_pointer == 125 && y_pointer == 53)
||(x_pointer == 126 && y_pointer == 53)
||(x_pointer == 127 && y_pointer == 53)
||(x_pointer == 128 && y_pointer == 53)
||(x_pointer == 129 && y_pointer == 53)
||(x_pointer == 130 && y_pointer == 53)
||(x_pointer == 29 && y_pointer == 54)
||(x_pointer == 30 && y_pointer == 54)
||(x_pointer == 31 && y_pointer == 54)
||(x_pointer == 32 && y_pointer == 54)
||(x_pointer == 33 && y_pointer == 54)
||(x_pointer == 34 && y_pointer == 54)
||(x_pointer == 35 && y_pointer == 54)
||(x_pointer == 36 && y_pointer == 54)
||(x_pointer == 37 && y_pointer == 54)
||(x_pointer == 38 && y_pointer == 54)
||(x_pointer == 39 && y_pointer == 54)
||(x_pointer == 40 && y_pointer == 54)
||(x_pointer == 41 && y_pointer == 54)
||(x_pointer == 42 && y_pointer == 54)
||(x_pointer == 43 && y_pointer == 54)
||(x_pointer == 44 && y_pointer == 54)
||(x_pointer == 45 && y_pointer == 54)
||(x_pointer == 46 && y_pointer == 54)
||(x_pointer == 47 && y_pointer == 54)
||(x_pointer == 48 && y_pointer == 54)
||(x_pointer == 49 && y_pointer == 54)
||(x_pointer == 50 && y_pointer == 54)
||(x_pointer == 51 && y_pointer == 54)
||(x_pointer == 52 && y_pointer == 54)
||(x_pointer == 53 && y_pointer == 54)
||(x_pointer == 54 && y_pointer == 54)
||(x_pointer == 55 && y_pointer == 54)
||(x_pointer == 56 && y_pointer == 54)
||(x_pointer == 57 && y_pointer == 54)
||(x_pointer == 58 && y_pointer == 54)
||(x_pointer == 59 && y_pointer == 54)
||(x_pointer == 60 && y_pointer == 54)
||(x_pointer == 61 && y_pointer == 54)
||(x_pointer == 62 && y_pointer == 54)
||(x_pointer == 63 && y_pointer == 54)
||(x_pointer == 64 && y_pointer == 54)
||(x_pointer == 65 && y_pointer == 54)
||(x_pointer == 66 && y_pointer == 54)
||(x_pointer == 67 && y_pointer == 54)
||(x_pointer == 92 && y_pointer == 54)
||(x_pointer == 93 && y_pointer == 54)
||(x_pointer == 94 && y_pointer == 54)
||(x_pointer == 95 && y_pointer == 54)
||(x_pointer == 96 && y_pointer == 54)
||(x_pointer == 97 && y_pointer == 54)
||(x_pointer == 98 && y_pointer == 54)
||(x_pointer == 99 && y_pointer == 54)
||(x_pointer == 100 && y_pointer == 54)
||(x_pointer == 101 && y_pointer == 54)
||(x_pointer == 102 && y_pointer == 54)
||(x_pointer == 103 && y_pointer == 54)
||(x_pointer == 104 && y_pointer == 54)
||(x_pointer == 105 && y_pointer == 54)
||(x_pointer == 106 && y_pointer == 54)
||(x_pointer == 107 && y_pointer == 54)
||(x_pointer == 108 && y_pointer == 54)
||(x_pointer == 109 && y_pointer == 54)
||(x_pointer == 110 && y_pointer == 54)
||(x_pointer == 111 && y_pointer == 54)
||(x_pointer == 112 && y_pointer == 54)
||(x_pointer == 113 && y_pointer == 54)
||(x_pointer == 114 && y_pointer == 54)
||(x_pointer == 115 && y_pointer == 54)
||(x_pointer == 116 && y_pointer == 54)
||(x_pointer == 117 && y_pointer == 54)
||(x_pointer == 118 && y_pointer == 54)
||(x_pointer == 119 && y_pointer == 54)
||(x_pointer == 120 && y_pointer == 54)
||(x_pointer == 121 && y_pointer == 54)
||(x_pointer == 122 && y_pointer == 54)
||(x_pointer == 123 && y_pointer == 54)
||(x_pointer == 124 && y_pointer == 54)
||(x_pointer == 125 && y_pointer == 54)
||(x_pointer == 126 && y_pointer == 54)
||(x_pointer == 127 && y_pointer == 54)
||(x_pointer == 128 && y_pointer == 54)
||(x_pointer == 129 && y_pointer == 54)
||(x_pointer == 130 && y_pointer == 54)
||(x_pointer == 29 && y_pointer == 55)
||(x_pointer == 30 && y_pointer == 55)
||(x_pointer == 31 && y_pointer == 55)
||(x_pointer == 32 && y_pointer == 55)
||(x_pointer == 33 && y_pointer == 55)
||(x_pointer == 34 && y_pointer == 55)
||(x_pointer == 35 && y_pointer == 55)
||(x_pointer == 36 && y_pointer == 55)
||(x_pointer == 37 && y_pointer == 55)
||(x_pointer == 38 && y_pointer == 55)
||(x_pointer == 39 && y_pointer == 55)
||(x_pointer == 40 && y_pointer == 55)
||(x_pointer == 41 && y_pointer == 55)
||(x_pointer == 42 && y_pointer == 55)
||(x_pointer == 43 && y_pointer == 55)
||(x_pointer == 44 && y_pointer == 55)
||(x_pointer == 45 && y_pointer == 55)
||(x_pointer == 46 && y_pointer == 55)
||(x_pointer == 47 && y_pointer == 55)
||(x_pointer == 48 && y_pointer == 55)
||(x_pointer == 49 && y_pointer == 55)
||(x_pointer == 50 && y_pointer == 55)
||(x_pointer == 51 && y_pointer == 55)
||(x_pointer == 52 && y_pointer == 55)
||(x_pointer == 53 && y_pointer == 55)
||(x_pointer == 54 && y_pointer == 55)
||(x_pointer == 55 && y_pointer == 55)
||(x_pointer == 56 && y_pointer == 55)
||(x_pointer == 57 && y_pointer == 55)
||(x_pointer == 58 && y_pointer == 55)
||(x_pointer == 59 && y_pointer == 55)
||(x_pointer == 60 && y_pointer == 55)
||(x_pointer == 61 && y_pointer == 55)
||(x_pointer == 62 && y_pointer == 55)
||(x_pointer == 63 && y_pointer == 55)
||(x_pointer == 64 && y_pointer == 55)
||(x_pointer == 65 && y_pointer == 55)
||(x_pointer == 66 && y_pointer == 55)
||(x_pointer == 67 && y_pointer == 55)
||(x_pointer == 92 && y_pointer == 55)
||(x_pointer == 93 && y_pointer == 55)
||(x_pointer == 94 && y_pointer == 55)
||(x_pointer == 95 && y_pointer == 55)
||(x_pointer == 96 && y_pointer == 55)
||(x_pointer == 97 && y_pointer == 55)
||(x_pointer == 98 && y_pointer == 55)
||(x_pointer == 99 && y_pointer == 55)
||(x_pointer == 100 && y_pointer == 55)
||(x_pointer == 101 && y_pointer == 55)
||(x_pointer == 102 && y_pointer == 55)
||(x_pointer == 103 && y_pointer == 55)
||(x_pointer == 104 && y_pointer == 55)
||(x_pointer == 105 && y_pointer == 55)
||(x_pointer == 106 && y_pointer == 55)
||(x_pointer == 107 && y_pointer == 55)
||(x_pointer == 108 && y_pointer == 55)
||(x_pointer == 109 && y_pointer == 55)
||(x_pointer == 110 && y_pointer == 55)
||(x_pointer == 111 && y_pointer == 55)
||(x_pointer == 112 && y_pointer == 55)
||(x_pointer == 113 && y_pointer == 55)
||(x_pointer == 114 && y_pointer == 55)
||(x_pointer == 115 && y_pointer == 55)
||(x_pointer == 116 && y_pointer == 55)
||(x_pointer == 117 && y_pointer == 55)
||(x_pointer == 118 && y_pointer == 55)
||(x_pointer == 119 && y_pointer == 55)
||(x_pointer == 120 && y_pointer == 55)
||(x_pointer == 121 && y_pointer == 55)
||(x_pointer == 122 && y_pointer == 55)
||(x_pointer == 123 && y_pointer == 55)
||(x_pointer == 124 && y_pointer == 55)
||(x_pointer == 125 && y_pointer == 55)
||(x_pointer == 126 && y_pointer == 55)
||(x_pointer == 127 && y_pointer == 55)
||(x_pointer == 128 && y_pointer == 55)
||(x_pointer == 129 && y_pointer == 55)
||(x_pointer == 130 && y_pointer == 55)
||(x_pointer == 29 && y_pointer == 56)
||(x_pointer == 30 && y_pointer == 56)
||(x_pointer == 31 && y_pointer == 56)
||(x_pointer == 32 && y_pointer == 56)
||(x_pointer == 33 && y_pointer == 56)
||(x_pointer == 34 && y_pointer == 56)
||(x_pointer == 35 && y_pointer == 56)
||(x_pointer == 36 && y_pointer == 56)
||(x_pointer == 37 && y_pointer == 56)
||(x_pointer == 38 && y_pointer == 56)
||(x_pointer == 39 && y_pointer == 56)
||(x_pointer == 40 && y_pointer == 56)
||(x_pointer == 41 && y_pointer == 56)
||(x_pointer == 42 && y_pointer == 56)
||(x_pointer == 43 && y_pointer == 56)
||(x_pointer == 44 && y_pointer == 56)
||(x_pointer == 45 && y_pointer == 56)
||(x_pointer == 46 && y_pointer == 56)
||(x_pointer == 47 && y_pointer == 56)
||(x_pointer == 48 && y_pointer == 56)
||(x_pointer == 49 && y_pointer == 56)
||(x_pointer == 50 && y_pointer == 56)
||(x_pointer == 51 && y_pointer == 56)
||(x_pointer == 52 && y_pointer == 56)
||(x_pointer == 53 && y_pointer == 56)
||(x_pointer == 54 && y_pointer == 56)
||(x_pointer == 55 && y_pointer == 56)
||(x_pointer == 56 && y_pointer == 56)
||(x_pointer == 57 && y_pointer == 56)
||(x_pointer == 58 && y_pointer == 56)
||(x_pointer == 59 && y_pointer == 56)
||(x_pointer == 60 && y_pointer == 56)
||(x_pointer == 61 && y_pointer == 56)
||(x_pointer == 62 && y_pointer == 56)
||(x_pointer == 63 && y_pointer == 56)
||(x_pointer == 64 && y_pointer == 56)
||(x_pointer == 65 && y_pointer == 56)
||(x_pointer == 66 && y_pointer == 56)
||(x_pointer == 67 && y_pointer == 56)
||(x_pointer == 92 && y_pointer == 56)
||(x_pointer == 93 && y_pointer == 56)
||(x_pointer == 94 && y_pointer == 56)
||(x_pointer == 95 && y_pointer == 56)
||(x_pointer == 96 && y_pointer == 56)
||(x_pointer == 97 && y_pointer == 56)
||(x_pointer == 98 && y_pointer == 56)
||(x_pointer == 99 && y_pointer == 56)
||(x_pointer == 100 && y_pointer == 56)
||(x_pointer == 101 && y_pointer == 56)
||(x_pointer == 102 && y_pointer == 56)
||(x_pointer == 103 && y_pointer == 56)
||(x_pointer == 104 && y_pointer == 56)
||(x_pointer == 105 && y_pointer == 56)
||(x_pointer == 106 && y_pointer == 56)
||(x_pointer == 107 && y_pointer == 56)
||(x_pointer == 108 && y_pointer == 56)
||(x_pointer == 109 && y_pointer == 56)
||(x_pointer == 110 && y_pointer == 56)
||(x_pointer == 111 && y_pointer == 56)
||(x_pointer == 112 && y_pointer == 56)
||(x_pointer == 113 && y_pointer == 56)
||(x_pointer == 114 && y_pointer == 56)
||(x_pointer == 115 && y_pointer == 56)
||(x_pointer == 116 && y_pointer == 56)
||(x_pointer == 117 && y_pointer == 56)
||(x_pointer == 118 && y_pointer == 56)
||(x_pointer == 119 && y_pointer == 56)
||(x_pointer == 120 && y_pointer == 56)
||(x_pointer == 121 && y_pointer == 56)
||(x_pointer == 122 && y_pointer == 56)
||(x_pointer == 123 && y_pointer == 56)
||(x_pointer == 124 && y_pointer == 56)
||(x_pointer == 125 && y_pointer == 56)
||(x_pointer == 126 && y_pointer == 56)
||(x_pointer == 127 && y_pointer == 56)
||(x_pointer == 128 && y_pointer == 56)
||(x_pointer == 129 && y_pointer == 56)
||(x_pointer == 130 && y_pointer == 56)
||(x_pointer == 29 && y_pointer == 57)
||(x_pointer == 30 && y_pointer == 57)
||(x_pointer == 31 && y_pointer == 57)
||(x_pointer == 32 && y_pointer == 57)
||(x_pointer == 33 && y_pointer == 57)
||(x_pointer == 34 && y_pointer == 57)
||(x_pointer == 35 && y_pointer == 57)
||(x_pointer == 36 && y_pointer == 57)
||(x_pointer == 37 && y_pointer == 57)
||(x_pointer == 38 && y_pointer == 57)
||(x_pointer == 39 && y_pointer == 57)
||(x_pointer == 40 && y_pointer == 57)
||(x_pointer == 41 && y_pointer == 57)
||(x_pointer == 42 && y_pointer == 57)
||(x_pointer == 43 && y_pointer == 57)
||(x_pointer == 44 && y_pointer == 57)
||(x_pointer == 45 && y_pointer == 57)
||(x_pointer == 46 && y_pointer == 57)
||(x_pointer == 47 && y_pointer == 57)
||(x_pointer == 48 && y_pointer == 57)
||(x_pointer == 49 && y_pointer == 57)
||(x_pointer == 50 && y_pointer == 57)
||(x_pointer == 51 && y_pointer == 57)
||(x_pointer == 52 && y_pointer == 57)
||(x_pointer == 53 && y_pointer == 57)
||(x_pointer == 54 && y_pointer == 57)
||(x_pointer == 55 && y_pointer == 57)
||(x_pointer == 56 && y_pointer == 57)
||(x_pointer == 57 && y_pointer == 57)
||(x_pointer == 58 && y_pointer == 57)
||(x_pointer == 59 && y_pointer == 57)
||(x_pointer == 60 && y_pointer == 57)
||(x_pointer == 61 && y_pointer == 57)
||(x_pointer == 62 && y_pointer == 57)
||(x_pointer == 63 && y_pointer == 57)
||(x_pointer == 64 && y_pointer == 57)
||(x_pointer == 65 && y_pointer == 57)
||(x_pointer == 66 && y_pointer == 57)
||(x_pointer == 67 && y_pointer == 57)
||(x_pointer == 92 && y_pointer == 57)
||(x_pointer == 93 && y_pointer == 57)
||(x_pointer == 94 && y_pointer == 57)
||(x_pointer == 95 && y_pointer == 57)
||(x_pointer == 96 && y_pointer == 57)
||(x_pointer == 97 && y_pointer == 57)
||(x_pointer == 98 && y_pointer == 57)
||(x_pointer == 99 && y_pointer == 57)
||(x_pointer == 100 && y_pointer == 57)
||(x_pointer == 101 && y_pointer == 57)
||(x_pointer == 102 && y_pointer == 57)
||(x_pointer == 103 && y_pointer == 57)
||(x_pointer == 104 && y_pointer == 57)
||(x_pointer == 105 && y_pointer == 57)
||(x_pointer == 106 && y_pointer == 57)
||(x_pointer == 107 && y_pointer == 57)
||(x_pointer == 108 && y_pointer == 57)
||(x_pointer == 109 && y_pointer == 57)
||(x_pointer == 110 && y_pointer == 57)
||(x_pointer == 111 && y_pointer == 57)
||(x_pointer == 112 && y_pointer == 57)
||(x_pointer == 113 && y_pointer == 57)
||(x_pointer == 114 && y_pointer == 57)
||(x_pointer == 115 && y_pointer == 57)
||(x_pointer == 116 && y_pointer == 57)
||(x_pointer == 117 && y_pointer == 57)
||(x_pointer == 118 && y_pointer == 57)
||(x_pointer == 119 && y_pointer == 57)
||(x_pointer == 120 && y_pointer == 57)
||(x_pointer == 121 && y_pointer == 57)
||(x_pointer == 122 && y_pointer == 57)
||(x_pointer == 123 && y_pointer == 57)
||(x_pointer == 124 && y_pointer == 57)
||(x_pointer == 125 && y_pointer == 57)
||(x_pointer == 126 && y_pointer == 57)
||(x_pointer == 127 && y_pointer == 57)
||(x_pointer == 128 && y_pointer == 57)
||(x_pointer == 129 && y_pointer == 57)
||(x_pointer == 130 && y_pointer == 57)
||(x_pointer == 29 && y_pointer == 58)
||(x_pointer == 30 && y_pointer == 58)
||(x_pointer == 31 && y_pointer == 58)
||(x_pointer == 32 && y_pointer == 58)
||(x_pointer == 33 && y_pointer == 58)
||(x_pointer == 34 && y_pointer == 58)
||(x_pointer == 35 && y_pointer == 58)
||(x_pointer == 36 && y_pointer == 58)
||(x_pointer == 37 && y_pointer == 58)
||(x_pointer == 38 && y_pointer == 58)
||(x_pointer == 39 && y_pointer == 58)
||(x_pointer == 40 && y_pointer == 58)
||(x_pointer == 41 && y_pointer == 58)
||(x_pointer == 42 && y_pointer == 58)
||(x_pointer == 43 && y_pointer == 58)
||(x_pointer == 44 && y_pointer == 58)
||(x_pointer == 45 && y_pointer == 58)
||(x_pointer == 46 && y_pointer == 58)
||(x_pointer == 47 && y_pointer == 58)
||(x_pointer == 48 && y_pointer == 58)
||(x_pointer == 49 && y_pointer == 58)
||(x_pointer == 50 && y_pointer == 58)
||(x_pointer == 51 && y_pointer == 58)
||(x_pointer == 52 && y_pointer == 58)
||(x_pointer == 53 && y_pointer == 58)
||(x_pointer == 54 && y_pointer == 58)
||(x_pointer == 55 && y_pointer == 58)
||(x_pointer == 56 && y_pointer == 58)
||(x_pointer == 57 && y_pointer == 58)
||(x_pointer == 58 && y_pointer == 58)
||(x_pointer == 59 && y_pointer == 58)
||(x_pointer == 60 && y_pointer == 58)
||(x_pointer == 61 && y_pointer == 58)
||(x_pointer == 62 && y_pointer == 58)
||(x_pointer == 63 && y_pointer == 58)
||(x_pointer == 64 && y_pointer == 58)
||(x_pointer == 65 && y_pointer == 58)
||(x_pointer == 66 && y_pointer == 58)
||(x_pointer == 67 && y_pointer == 58)
||(x_pointer == 92 && y_pointer == 58)
||(x_pointer == 93 && y_pointer == 58)
||(x_pointer == 94 && y_pointer == 58)
||(x_pointer == 95 && y_pointer == 58)
||(x_pointer == 96 && y_pointer == 58)
||(x_pointer == 97 && y_pointer == 58)
||(x_pointer == 98 && y_pointer == 58)
||(x_pointer == 99 && y_pointer == 58)
||(x_pointer == 100 && y_pointer == 58)
||(x_pointer == 101 && y_pointer == 58)
||(x_pointer == 102 && y_pointer == 58)
||(x_pointer == 103 && y_pointer == 58)
||(x_pointer == 104 && y_pointer == 58)
||(x_pointer == 105 && y_pointer == 58)
||(x_pointer == 106 && y_pointer == 58)
||(x_pointer == 107 && y_pointer == 58)
||(x_pointer == 108 && y_pointer == 58)
||(x_pointer == 109 && y_pointer == 58)
||(x_pointer == 110 && y_pointer == 58)
||(x_pointer == 111 && y_pointer == 58)
||(x_pointer == 112 && y_pointer == 58)
||(x_pointer == 113 && y_pointer == 58)
||(x_pointer == 114 && y_pointer == 58)
||(x_pointer == 115 && y_pointer == 58)
||(x_pointer == 116 && y_pointer == 58)
||(x_pointer == 117 && y_pointer == 58)
||(x_pointer == 118 && y_pointer == 58)
||(x_pointer == 119 && y_pointer == 58)
||(x_pointer == 120 && y_pointer == 58)
||(x_pointer == 121 && y_pointer == 58)
||(x_pointer == 122 && y_pointer == 58)
||(x_pointer == 123 && y_pointer == 58)
||(x_pointer == 124 && y_pointer == 58)
||(x_pointer == 125 && y_pointer == 58)
||(x_pointer == 126 && y_pointer == 58)
||(x_pointer == 127 && y_pointer == 58)
||(x_pointer == 128 && y_pointer == 58)
||(x_pointer == 129 && y_pointer == 58)
||(x_pointer == 130 && y_pointer == 58));
	wire barrier_pixel_2 = current_level == 2 && ((x_pointer == 2 && y_pointer == 2)
||(x_pointer == 3 && y_pointer == 2)
||(x_pointer == 4 && y_pointer == 2)
||(x_pointer == 5 && y_pointer == 2)
||(x_pointer == 6 && y_pointer == 2)
||(x_pointer == 7 && y_pointer == 2)
||(x_pointer == 8 && y_pointer == 2)
||(x_pointer == 9 && y_pointer == 2)
||(x_pointer == 10 && y_pointer == 2)
||(x_pointer == 11 && y_pointer == 2)
||(x_pointer == 12 && y_pointer == 2)
||(x_pointer == 13 && y_pointer == 2)
||(x_pointer == 14 && y_pointer == 2)
||(x_pointer == 15 && y_pointer == 2)
||(x_pointer == 16 && y_pointer == 2)
||(x_pointer == 17 && y_pointer == 2)
||(x_pointer == 18 && y_pointer == 2)
||(x_pointer == 19 && y_pointer == 2)
||(x_pointer == 20 && y_pointer == 2)
||(x_pointer == 21 && y_pointer == 2)
||(x_pointer == 22 && y_pointer == 2)
||(x_pointer == 23 && y_pointer == 2)
||(x_pointer == 24 && y_pointer == 2)
||(x_pointer == 25 && y_pointer == 2)
||(x_pointer == 26 && y_pointer == 2)
||(x_pointer == 27 && y_pointer == 2)
||(x_pointer == 28 && y_pointer == 2)
||(x_pointer == 29 && y_pointer == 2)
||(x_pointer == 30 && y_pointer == 2)
||(x_pointer == 31 && y_pointer == 2)
||(x_pointer == 32 && y_pointer == 2)
||(x_pointer == 33 && y_pointer == 2)
||(x_pointer == 34 && y_pointer == 2)
||(x_pointer == 35 && y_pointer == 2)
||(x_pointer == 36 && y_pointer == 2)
||(x_pointer == 37 && y_pointer == 2)
||(x_pointer == 38 && y_pointer == 2)
||(x_pointer == 39 && y_pointer == 2)
||(x_pointer == 40 && y_pointer == 2)
||(x_pointer == 41 && y_pointer == 2)
||(x_pointer == 42 && y_pointer == 2)
||(x_pointer == 43 && y_pointer == 2)
||(x_pointer == 44 && y_pointer == 2)
||(x_pointer == 45 && y_pointer == 2)
||(x_pointer == 46 && y_pointer == 2)
||(x_pointer == 47 && y_pointer == 2)
||(x_pointer == 48 && y_pointer == 2)
||(x_pointer == 49 && y_pointer == 2)
||(x_pointer == 50 && y_pointer == 2)
||(x_pointer == 51 && y_pointer == 2)
||(x_pointer == 52 && y_pointer == 2)
||(x_pointer == 53 && y_pointer == 2)
||(x_pointer == 54 && y_pointer == 2)
||(x_pointer == 55 && y_pointer == 2)
||(x_pointer == 56 && y_pointer == 2)
||(x_pointer == 57 && y_pointer == 2)
||(x_pointer == 58 && y_pointer == 2)
||(x_pointer == 59 && y_pointer == 2)
||(x_pointer == 60 && y_pointer == 2)
||(x_pointer == 61 && y_pointer == 2)
||(x_pointer == 62 && y_pointer == 2)
||(x_pointer == 63 && y_pointer == 2)
||(x_pointer == 64 && y_pointer == 2)
||(x_pointer == 65 && y_pointer == 2)
||(x_pointer == 66 && y_pointer == 2)
||(x_pointer == 67 && y_pointer == 2)
||(x_pointer == 68 && y_pointer == 2)
||(x_pointer == 69 && y_pointer == 2)
||(x_pointer == 70 && y_pointer == 2)
||(x_pointer == 71 && y_pointer == 2)
||(x_pointer == 72 && y_pointer == 2)
||(x_pointer == 73 && y_pointer == 2)
||(x_pointer == 74 && y_pointer == 2)
||(x_pointer == 75 && y_pointer == 2)
||(x_pointer == 76 && y_pointer == 2)
||(x_pointer == 77 && y_pointer == 2)
||(x_pointer == 78 && y_pointer == 2)
||(x_pointer == 79 && y_pointer == 2)
||(x_pointer == 80 && y_pointer == 2)
||(x_pointer == 81 && y_pointer == 2)
||(x_pointer == 82 && y_pointer == 2)
||(x_pointer == 83 && y_pointer == 2)
||(x_pointer == 84 && y_pointer == 2)
||(x_pointer == 85 && y_pointer == 2)
||(x_pointer == 86 && y_pointer == 2)
||(x_pointer == 87 && y_pointer == 2)
||(x_pointer == 88 && y_pointer == 2)
||(x_pointer == 89 && y_pointer == 2)
||(x_pointer == 90 && y_pointer == 2)
||(x_pointer == 91 && y_pointer == 2)
||(x_pointer == 92 && y_pointer == 2)
||(x_pointer == 93 && y_pointer == 2)
||(x_pointer == 94 && y_pointer == 2)
||(x_pointer == 95 && y_pointer == 2)
||(x_pointer == 96 && y_pointer == 2)
||(x_pointer == 97 && y_pointer == 2)
||(x_pointer == 98 && y_pointer == 2)
||(x_pointer == 99 && y_pointer == 2)
||(x_pointer == 100 && y_pointer == 2)
||(x_pointer == 101 && y_pointer == 2)
||(x_pointer == 102 && y_pointer == 2)
||(x_pointer == 103 && y_pointer == 2)
||(x_pointer == 104 && y_pointer == 2)
||(x_pointer == 105 && y_pointer == 2)
||(x_pointer == 106 && y_pointer == 2)
||(x_pointer == 107 && y_pointer == 2)
||(x_pointer == 108 && y_pointer == 2)
||(x_pointer == 109 && y_pointer == 2)
||(x_pointer == 110 && y_pointer == 2)
||(x_pointer == 111 && y_pointer == 2)
||(x_pointer == 112 && y_pointer == 2)
||(x_pointer == 113 && y_pointer == 2)
||(x_pointer == 114 && y_pointer == 2)
||(x_pointer == 115 && y_pointer == 2)
||(x_pointer == 116 && y_pointer == 2)
||(x_pointer == 117 && y_pointer == 2)
||(x_pointer == 118 && y_pointer == 2)
||(x_pointer == 119 && y_pointer == 2)
||(x_pointer == 120 && y_pointer == 2)
||(x_pointer == 121 && y_pointer == 2)
||(x_pointer == 122 && y_pointer == 2)
||(x_pointer == 123 && y_pointer == 2)
||(x_pointer == 124 && y_pointer == 2)
||(x_pointer == 125 && y_pointer == 2)
||(x_pointer == 126 && y_pointer == 2)
||(x_pointer == 127 && y_pointer == 2)
||(x_pointer == 128 && y_pointer == 2)
||(x_pointer == 129 && y_pointer == 2)
||(x_pointer == 130 && y_pointer == 2)
||(x_pointer == 131 && y_pointer == 2)
||(x_pointer == 132 && y_pointer == 2)
||(x_pointer == 133 && y_pointer == 2)
||(x_pointer == 134 && y_pointer == 2)
||(x_pointer == 135 && y_pointer == 2)
||(x_pointer == 136 && y_pointer == 2)
||(x_pointer == 137 && y_pointer == 2)
||(x_pointer == 138 && y_pointer == 2)
||(x_pointer == 139 && y_pointer == 2)
||(x_pointer == 140 && y_pointer == 2)
||(x_pointer == 141 && y_pointer == 2)
||(x_pointer == 142 && y_pointer == 2)
||(x_pointer == 143 && y_pointer == 2)
||(x_pointer == 144 && y_pointer == 2)
||(x_pointer == 145 && y_pointer == 2)
||(x_pointer == 146 && y_pointer == 2)
||(x_pointer == 147 && y_pointer == 2)
||(x_pointer == 148 && y_pointer == 2)
||(x_pointer == 149 && y_pointer == 2)
||(x_pointer == 150 && y_pointer == 2)
||(x_pointer == 151 && y_pointer == 2)
||(x_pointer == 152 && y_pointer == 2)
||(x_pointer == 153 && y_pointer == 2)
||(x_pointer == 154 && y_pointer == 2)
||(x_pointer == 155 && y_pointer == 2)
||(x_pointer == 156 && y_pointer == 2)
||(x_pointer == 157 && y_pointer == 2)
||(x_pointer == 2 && y_pointer == 3)
||(x_pointer == 3 && y_pointer == 3)
||(x_pointer == 4 && y_pointer == 3)
||(x_pointer == 5 && y_pointer == 3)
||(x_pointer == 6 && y_pointer == 3)
||(x_pointer == 7 && y_pointer == 3)
||(x_pointer == 8 && y_pointer == 3)
||(x_pointer == 9 && y_pointer == 3)
||(x_pointer == 10 && y_pointer == 3)
||(x_pointer == 11 && y_pointer == 3)
||(x_pointer == 12 && y_pointer == 3)
||(x_pointer == 13 && y_pointer == 3)
||(x_pointer == 14 && y_pointer == 3)
||(x_pointer == 15 && y_pointer == 3)
||(x_pointer == 16 && y_pointer == 3)
||(x_pointer == 17 && y_pointer == 3)
||(x_pointer == 18 && y_pointer == 3)
||(x_pointer == 19 && y_pointer == 3)
||(x_pointer == 20 && y_pointer == 3)
||(x_pointer == 21 && y_pointer == 3)
||(x_pointer == 22 && y_pointer == 3)
||(x_pointer == 23 && y_pointer == 3)
||(x_pointer == 24 && y_pointer == 3)
||(x_pointer == 25 && y_pointer == 3)
||(x_pointer == 26 && y_pointer == 3)
||(x_pointer == 27 && y_pointer == 3)
||(x_pointer == 28 && y_pointer == 3)
||(x_pointer == 29 && y_pointer == 3)
||(x_pointer == 30 && y_pointer == 3)
||(x_pointer == 31 && y_pointer == 3)
||(x_pointer == 32 && y_pointer == 3)
||(x_pointer == 33 && y_pointer == 3)
||(x_pointer == 34 && y_pointer == 3)
||(x_pointer == 35 && y_pointer == 3)
||(x_pointer == 36 && y_pointer == 3)
||(x_pointer == 37 && y_pointer == 3)
||(x_pointer == 38 && y_pointer == 3)
||(x_pointer == 39 && y_pointer == 3)
||(x_pointer == 40 && y_pointer == 3)
||(x_pointer == 41 && y_pointer == 3)
||(x_pointer == 42 && y_pointer == 3)
||(x_pointer == 43 && y_pointer == 3)
||(x_pointer == 44 && y_pointer == 3)
||(x_pointer == 45 && y_pointer == 3)
||(x_pointer == 46 && y_pointer == 3)
||(x_pointer == 47 && y_pointer == 3)
||(x_pointer == 48 && y_pointer == 3)
||(x_pointer == 49 && y_pointer == 3)
||(x_pointer == 50 && y_pointer == 3)
||(x_pointer == 51 && y_pointer == 3)
||(x_pointer == 52 && y_pointer == 3)
||(x_pointer == 53 && y_pointer == 3)
||(x_pointer == 54 && y_pointer == 3)
||(x_pointer == 55 && y_pointer == 3)
||(x_pointer == 56 && y_pointer == 3)
||(x_pointer == 57 && y_pointer == 3)
||(x_pointer == 58 && y_pointer == 3)
||(x_pointer == 59 && y_pointer == 3)
||(x_pointer == 60 && y_pointer == 3)
||(x_pointer == 61 && y_pointer == 3)
||(x_pointer == 62 && y_pointer == 3)
||(x_pointer == 63 && y_pointer == 3)
||(x_pointer == 64 && y_pointer == 3)
||(x_pointer == 65 && y_pointer == 3)
||(x_pointer == 66 && y_pointer == 3)
||(x_pointer == 67 && y_pointer == 3)
||(x_pointer == 68 && y_pointer == 3)
||(x_pointer == 69 && y_pointer == 3)
||(x_pointer == 70 && y_pointer == 3)
||(x_pointer == 71 && y_pointer == 3)
||(x_pointer == 72 && y_pointer == 3)
||(x_pointer == 73 && y_pointer == 3)
||(x_pointer == 74 && y_pointer == 3)
||(x_pointer == 75 && y_pointer == 3)
||(x_pointer == 76 && y_pointer == 3)
||(x_pointer == 77 && y_pointer == 3)
||(x_pointer == 78 && y_pointer == 3)
||(x_pointer == 79 && y_pointer == 3)
||(x_pointer == 80 && y_pointer == 3)
||(x_pointer == 81 && y_pointer == 3)
||(x_pointer == 82 && y_pointer == 3)
||(x_pointer == 83 && y_pointer == 3)
||(x_pointer == 84 && y_pointer == 3)
||(x_pointer == 85 && y_pointer == 3)
||(x_pointer == 86 && y_pointer == 3)
||(x_pointer == 87 && y_pointer == 3)
||(x_pointer == 88 && y_pointer == 3)
||(x_pointer == 89 && y_pointer == 3)
||(x_pointer == 90 && y_pointer == 3)
||(x_pointer == 91 && y_pointer == 3)
||(x_pointer == 92 && y_pointer == 3)
||(x_pointer == 93 && y_pointer == 3)
||(x_pointer == 94 && y_pointer == 3)
||(x_pointer == 95 && y_pointer == 3)
||(x_pointer == 96 && y_pointer == 3)
||(x_pointer == 97 && y_pointer == 3)
||(x_pointer == 98 && y_pointer == 3)
||(x_pointer == 99 && y_pointer == 3)
||(x_pointer == 100 && y_pointer == 3)
||(x_pointer == 101 && y_pointer == 3)
||(x_pointer == 102 && y_pointer == 3)
||(x_pointer == 103 && y_pointer == 3)
||(x_pointer == 104 && y_pointer == 3)
||(x_pointer == 105 && y_pointer == 3)
||(x_pointer == 106 && y_pointer == 3)
||(x_pointer == 107 && y_pointer == 3)
||(x_pointer == 108 && y_pointer == 3)
||(x_pointer == 109 && y_pointer == 3)
||(x_pointer == 110 && y_pointer == 3)
||(x_pointer == 111 && y_pointer == 3)
||(x_pointer == 112 && y_pointer == 3)
||(x_pointer == 113 && y_pointer == 3)
||(x_pointer == 114 && y_pointer == 3)
||(x_pointer == 115 && y_pointer == 3)
||(x_pointer == 116 && y_pointer == 3)
||(x_pointer == 117 && y_pointer == 3)
||(x_pointer == 118 && y_pointer == 3)
||(x_pointer == 119 && y_pointer == 3)
||(x_pointer == 120 && y_pointer == 3)
||(x_pointer == 121 && y_pointer == 3)
||(x_pointer == 122 && y_pointer == 3)
||(x_pointer == 123 && y_pointer == 3)
||(x_pointer == 124 && y_pointer == 3)
||(x_pointer == 125 && y_pointer == 3)
||(x_pointer == 126 && y_pointer == 3)
||(x_pointer == 127 && y_pointer == 3)
||(x_pointer == 128 && y_pointer == 3)
||(x_pointer == 129 && y_pointer == 3)
||(x_pointer == 130 && y_pointer == 3)
||(x_pointer == 131 && y_pointer == 3)
||(x_pointer == 132 && y_pointer == 3)
||(x_pointer == 133 && y_pointer == 3)
||(x_pointer == 134 && y_pointer == 3)
||(x_pointer == 135 && y_pointer == 3)
||(x_pointer == 136 && y_pointer == 3)
||(x_pointer == 137 && y_pointer == 3)
||(x_pointer == 138 && y_pointer == 3)
||(x_pointer == 139 && y_pointer == 3)
||(x_pointer == 140 && y_pointer == 3)
||(x_pointer == 141 && y_pointer == 3)
||(x_pointer == 142 && y_pointer == 3)
||(x_pointer == 143 && y_pointer == 3)
||(x_pointer == 144 && y_pointer == 3)
||(x_pointer == 145 && y_pointer == 3)
||(x_pointer == 146 && y_pointer == 3)
||(x_pointer == 147 && y_pointer == 3)
||(x_pointer == 148 && y_pointer == 3)
||(x_pointer == 149 && y_pointer == 3)
||(x_pointer == 150 && y_pointer == 3)
||(x_pointer == 151 && y_pointer == 3)
||(x_pointer == 152 && y_pointer == 3)
||(x_pointer == 153 && y_pointer == 3)
||(x_pointer == 154 && y_pointer == 3)
||(x_pointer == 155 && y_pointer == 3)
||(x_pointer == 156 && y_pointer == 3)
||(x_pointer == 157 && y_pointer == 3)
||(x_pointer == 2 && y_pointer == 4)
||(x_pointer == 3 && y_pointer == 4)
||(x_pointer == 4 && y_pointer == 4)
||(x_pointer == 5 && y_pointer == 4)
||(x_pointer == 6 && y_pointer == 4)
||(x_pointer == 7 && y_pointer == 4)
||(x_pointer == 8 && y_pointer == 4)
||(x_pointer == 9 && y_pointer == 4)
||(x_pointer == 10 && y_pointer == 4)
||(x_pointer == 11 && y_pointer == 4)
||(x_pointer == 12 && y_pointer == 4)
||(x_pointer == 13 && y_pointer == 4)
||(x_pointer == 14 && y_pointer == 4)
||(x_pointer == 15 && y_pointer == 4)
||(x_pointer == 16 && y_pointer == 4)
||(x_pointer == 17 && y_pointer == 4)
||(x_pointer == 18 && y_pointer == 4)
||(x_pointer == 19 && y_pointer == 4)
||(x_pointer == 20 && y_pointer == 4)
||(x_pointer == 21 && y_pointer == 4)
||(x_pointer == 22 && y_pointer == 4)
||(x_pointer == 23 && y_pointer == 4)
||(x_pointer == 24 && y_pointer == 4)
||(x_pointer == 25 && y_pointer == 4)
||(x_pointer == 26 && y_pointer == 4)
||(x_pointer == 27 && y_pointer == 4)
||(x_pointer == 28 && y_pointer == 4)
||(x_pointer == 29 && y_pointer == 4)
||(x_pointer == 30 && y_pointer == 4)
||(x_pointer == 31 && y_pointer == 4)
||(x_pointer == 32 && y_pointer == 4)
||(x_pointer == 33 && y_pointer == 4)
||(x_pointer == 34 && y_pointer == 4)
||(x_pointer == 35 && y_pointer == 4)
||(x_pointer == 36 && y_pointer == 4)
||(x_pointer == 37 && y_pointer == 4)
||(x_pointer == 38 && y_pointer == 4)
||(x_pointer == 39 && y_pointer == 4)
||(x_pointer == 40 && y_pointer == 4)
||(x_pointer == 41 && y_pointer == 4)
||(x_pointer == 42 && y_pointer == 4)
||(x_pointer == 43 && y_pointer == 4)
||(x_pointer == 44 && y_pointer == 4)
||(x_pointer == 45 && y_pointer == 4)
||(x_pointer == 46 && y_pointer == 4)
||(x_pointer == 47 && y_pointer == 4)
||(x_pointer == 48 && y_pointer == 4)
||(x_pointer == 49 && y_pointer == 4)
||(x_pointer == 50 && y_pointer == 4)
||(x_pointer == 51 && y_pointer == 4)
||(x_pointer == 52 && y_pointer == 4)
||(x_pointer == 53 && y_pointer == 4)
||(x_pointer == 54 && y_pointer == 4)
||(x_pointer == 55 && y_pointer == 4)
||(x_pointer == 56 && y_pointer == 4)
||(x_pointer == 57 && y_pointer == 4)
||(x_pointer == 58 && y_pointer == 4)
||(x_pointer == 59 && y_pointer == 4)
||(x_pointer == 60 && y_pointer == 4)
||(x_pointer == 61 && y_pointer == 4)
||(x_pointer == 62 && y_pointer == 4)
||(x_pointer == 63 && y_pointer == 4)
||(x_pointer == 64 && y_pointer == 4)
||(x_pointer == 65 && y_pointer == 4)
||(x_pointer == 66 && y_pointer == 4)
||(x_pointer == 67 && y_pointer == 4)
||(x_pointer == 68 && y_pointer == 4)
||(x_pointer == 69 && y_pointer == 4)
||(x_pointer == 70 && y_pointer == 4)
||(x_pointer == 71 && y_pointer == 4)
||(x_pointer == 72 && y_pointer == 4)
||(x_pointer == 73 && y_pointer == 4)
||(x_pointer == 74 && y_pointer == 4)
||(x_pointer == 75 && y_pointer == 4)
||(x_pointer == 76 && y_pointer == 4)
||(x_pointer == 77 && y_pointer == 4)
||(x_pointer == 78 && y_pointer == 4)
||(x_pointer == 79 && y_pointer == 4)
||(x_pointer == 80 && y_pointer == 4)
||(x_pointer == 81 && y_pointer == 4)
||(x_pointer == 82 && y_pointer == 4)
||(x_pointer == 83 && y_pointer == 4)
||(x_pointer == 84 && y_pointer == 4)
||(x_pointer == 85 && y_pointer == 4)
||(x_pointer == 86 && y_pointer == 4)
||(x_pointer == 87 && y_pointer == 4)
||(x_pointer == 88 && y_pointer == 4)
||(x_pointer == 89 && y_pointer == 4)
||(x_pointer == 90 && y_pointer == 4)
||(x_pointer == 91 && y_pointer == 4)
||(x_pointer == 92 && y_pointer == 4)
||(x_pointer == 93 && y_pointer == 4)
||(x_pointer == 94 && y_pointer == 4)
||(x_pointer == 95 && y_pointer == 4)
||(x_pointer == 96 && y_pointer == 4)
||(x_pointer == 97 && y_pointer == 4)
||(x_pointer == 98 && y_pointer == 4)
||(x_pointer == 99 && y_pointer == 4)
||(x_pointer == 100 && y_pointer == 4)
||(x_pointer == 101 && y_pointer == 4)
||(x_pointer == 102 && y_pointer == 4)
||(x_pointer == 103 && y_pointer == 4)
||(x_pointer == 104 && y_pointer == 4)
||(x_pointer == 105 && y_pointer == 4)
||(x_pointer == 106 && y_pointer == 4)
||(x_pointer == 107 && y_pointer == 4)
||(x_pointer == 108 && y_pointer == 4)
||(x_pointer == 109 && y_pointer == 4)
||(x_pointer == 110 && y_pointer == 4)
||(x_pointer == 111 && y_pointer == 4)
||(x_pointer == 112 && y_pointer == 4)
||(x_pointer == 113 && y_pointer == 4)
||(x_pointer == 114 && y_pointer == 4)
||(x_pointer == 115 && y_pointer == 4)
||(x_pointer == 116 && y_pointer == 4)
||(x_pointer == 117 && y_pointer == 4)
||(x_pointer == 118 && y_pointer == 4)
||(x_pointer == 119 && y_pointer == 4)
||(x_pointer == 120 && y_pointer == 4)
||(x_pointer == 121 && y_pointer == 4)
||(x_pointer == 122 && y_pointer == 4)
||(x_pointer == 123 && y_pointer == 4)
||(x_pointer == 124 && y_pointer == 4)
||(x_pointer == 125 && y_pointer == 4)
||(x_pointer == 126 && y_pointer == 4)
||(x_pointer == 127 && y_pointer == 4)
||(x_pointer == 128 && y_pointer == 4)
||(x_pointer == 129 && y_pointer == 4)
||(x_pointer == 130 && y_pointer == 4)
||(x_pointer == 131 && y_pointer == 4)
||(x_pointer == 132 && y_pointer == 4)
||(x_pointer == 133 && y_pointer == 4)
||(x_pointer == 134 && y_pointer == 4)
||(x_pointer == 135 && y_pointer == 4)
||(x_pointer == 136 && y_pointer == 4)
||(x_pointer == 137 && y_pointer == 4)
||(x_pointer == 138 && y_pointer == 4)
||(x_pointer == 139 && y_pointer == 4)
||(x_pointer == 140 && y_pointer == 4)
||(x_pointer == 141 && y_pointer == 4)
||(x_pointer == 142 && y_pointer == 4)
||(x_pointer == 143 && y_pointer == 4)
||(x_pointer == 144 && y_pointer == 4)
||(x_pointer == 145 && y_pointer == 4)
||(x_pointer == 146 && y_pointer == 4)
||(x_pointer == 147 && y_pointer == 4)
||(x_pointer == 148 && y_pointer == 4)
||(x_pointer == 149 && y_pointer == 4)
||(x_pointer == 150 && y_pointer == 4)
||(x_pointer == 151 && y_pointer == 4)
||(x_pointer == 152 && y_pointer == 4)
||(x_pointer == 153 && y_pointer == 4)
||(x_pointer == 154 && y_pointer == 4)
||(x_pointer == 155 && y_pointer == 4)
||(x_pointer == 156 && y_pointer == 4)
||(x_pointer == 157 && y_pointer == 4)
||(x_pointer == 2 && y_pointer == 5)
||(x_pointer == 3 && y_pointer == 5)
||(x_pointer == 4 && y_pointer == 5)
||(x_pointer == 155 && y_pointer == 5)
||(x_pointer == 156 && y_pointer == 5)
||(x_pointer == 157 && y_pointer == 5)
||(x_pointer == 2 && y_pointer == 6)
||(x_pointer == 3 && y_pointer == 6)
||(x_pointer == 4 && y_pointer == 6)
||(x_pointer == 155 && y_pointer == 6)
||(x_pointer == 156 && y_pointer == 6)
||(x_pointer == 157 && y_pointer == 6)
||(x_pointer == 2 && y_pointer == 7)
||(x_pointer == 3 && y_pointer == 7)
||(x_pointer == 4 && y_pointer == 7)
||(x_pointer == 155 && y_pointer == 7)
||(x_pointer == 156 && y_pointer == 7)
||(x_pointer == 157 && y_pointer == 7)
||(x_pointer == 2 && y_pointer == 8)
||(x_pointer == 3 && y_pointer == 8)
||(x_pointer == 4 && y_pointer == 8)
||(x_pointer == 155 && y_pointer == 8)
||(x_pointer == 156 && y_pointer == 8)
||(x_pointer == 157 && y_pointer == 8)
||(x_pointer == 2 && y_pointer == 9)
||(x_pointer == 3 && y_pointer == 9)
||(x_pointer == 4 && y_pointer == 9)
||(x_pointer == 155 && y_pointer == 9)
||(x_pointer == 156 && y_pointer == 9)
||(x_pointer == 157 && y_pointer == 9)
||(x_pointer == 2 && y_pointer == 10)
||(x_pointer == 3 && y_pointer == 10)
||(x_pointer == 4 && y_pointer == 10)
||(x_pointer == 155 && y_pointer == 10)
||(x_pointer == 156 && y_pointer == 10)
||(x_pointer == 157 && y_pointer == 10)
||(x_pointer == 2 && y_pointer == 11)
||(x_pointer == 3 && y_pointer == 11)
||(x_pointer == 4 && y_pointer == 11)
||(x_pointer == 155 && y_pointer == 11)
||(x_pointer == 156 && y_pointer == 11)
||(x_pointer == 157 && y_pointer == 11)
||(x_pointer == 2 && y_pointer == 12)
||(x_pointer == 3 && y_pointer == 12)
||(x_pointer == 4 && y_pointer == 12)
||(x_pointer == 155 && y_pointer == 12)
||(x_pointer == 156 && y_pointer == 12)
||(x_pointer == 157 && y_pointer == 12)
||(x_pointer == 2 && y_pointer == 13)
||(x_pointer == 3 && y_pointer == 13)
||(x_pointer == 4 && y_pointer == 13)
||(x_pointer == 155 && y_pointer == 13)
||(x_pointer == 156 && y_pointer == 13)
||(x_pointer == 157 && y_pointer == 13)
||(x_pointer == 2 && y_pointer == 14)
||(x_pointer == 3 && y_pointer == 14)
||(x_pointer == 4 && y_pointer == 14)
||(x_pointer == 155 && y_pointer == 14)
||(x_pointer == 156 && y_pointer == 14)
||(x_pointer == 157 && y_pointer == 14)
||(x_pointer == 2 && y_pointer == 15)
||(x_pointer == 3 && y_pointer == 15)
||(x_pointer == 4 && y_pointer == 15)
||(x_pointer == 155 && y_pointer == 15)
||(x_pointer == 156 && y_pointer == 15)
||(x_pointer == 157 && y_pointer == 15)
||(x_pointer == 2 && y_pointer == 16)
||(x_pointer == 3 && y_pointer == 16)
||(x_pointer == 4 && y_pointer == 16)
||(x_pointer == 155 && y_pointer == 16)
||(x_pointer == 156 && y_pointer == 16)
||(x_pointer == 157 && y_pointer == 16)
||(x_pointer == 2 && y_pointer == 17)
||(x_pointer == 3 && y_pointer == 17)
||(x_pointer == 4 && y_pointer == 17)
||(x_pointer == 155 && y_pointer == 17)
||(x_pointer == 156 && y_pointer == 17)
||(x_pointer == 157 && y_pointer == 17)
||(x_pointer == 2 && y_pointer == 18)
||(x_pointer == 3 && y_pointer == 18)
||(x_pointer == 4 && y_pointer == 18)
||(x_pointer == 155 && y_pointer == 18)
||(x_pointer == 156 && y_pointer == 18)
||(x_pointer == 157 && y_pointer == 18)
||(x_pointer == 2 && y_pointer == 19)
||(x_pointer == 3 && y_pointer == 19)
||(x_pointer == 4 && y_pointer == 19)
||(x_pointer == 155 && y_pointer == 19)
||(x_pointer == 156 && y_pointer == 19)
||(x_pointer == 157 && y_pointer == 19)
||(x_pointer == 2 && y_pointer == 20)
||(x_pointer == 3 && y_pointer == 20)
||(x_pointer == 4 && y_pointer == 20)
||(x_pointer == 155 && y_pointer == 20)
||(x_pointer == 156 && y_pointer == 20)
||(x_pointer == 157 && y_pointer == 20)
||(x_pointer == 2 && y_pointer == 21)
||(x_pointer == 3 && y_pointer == 21)
||(x_pointer == 4 && y_pointer == 21)
||(x_pointer == 155 && y_pointer == 21)
||(x_pointer == 156 && y_pointer == 21)
||(x_pointer == 157 && y_pointer == 21)
||(x_pointer == 2 && y_pointer == 22)
||(x_pointer == 3 && y_pointer == 22)
||(x_pointer == 4 && y_pointer == 22)
||(x_pointer == 155 && y_pointer == 22)
||(x_pointer == 156 && y_pointer == 22)
||(x_pointer == 157 && y_pointer == 22)
||(x_pointer == 2 && y_pointer == 23)
||(x_pointer == 3 && y_pointer == 23)
||(x_pointer == 4 && y_pointer == 23)
||(x_pointer == 50 && y_pointer == 23)
||(x_pointer == 51 && y_pointer == 23)
||(x_pointer == 52 && y_pointer == 23)
||(x_pointer == 53 && y_pointer == 23)
||(x_pointer == 54 && y_pointer == 23)
||(x_pointer == 55 && y_pointer == 23)
||(x_pointer == 56 && y_pointer == 23)
||(x_pointer == 57 && y_pointer == 23)
||(x_pointer == 58 && y_pointer == 23)
||(x_pointer == 59 && y_pointer == 23)
||(x_pointer == 60 && y_pointer == 23)
||(x_pointer == 61 && y_pointer == 23)
||(x_pointer == 62 && y_pointer == 23)
||(x_pointer == 63 && y_pointer == 23)
||(x_pointer == 64 && y_pointer == 23)
||(x_pointer == 65 && y_pointer == 23)
||(x_pointer == 66 && y_pointer == 23)
||(x_pointer == 67 && y_pointer == 23)
||(x_pointer == 68 && y_pointer == 23)
||(x_pointer == 69 && y_pointer == 23)
||(x_pointer == 70 && y_pointer == 23)
||(x_pointer == 71 && y_pointer == 23)
||(x_pointer == 72 && y_pointer == 23)
||(x_pointer == 73 && y_pointer == 23)
||(x_pointer == 89 && y_pointer == 23)
||(x_pointer == 90 && y_pointer == 23)
||(x_pointer == 91 && y_pointer == 23)
||(x_pointer == 92 && y_pointer == 23)
||(x_pointer == 93 && y_pointer == 23)
||(x_pointer == 94 && y_pointer == 23)
||(x_pointer == 95 && y_pointer == 23)
||(x_pointer == 96 && y_pointer == 23)
||(x_pointer == 97 && y_pointer == 23)
||(x_pointer == 98 && y_pointer == 23)
||(x_pointer == 99 && y_pointer == 23)
||(x_pointer == 100 && y_pointer == 23)
||(x_pointer == 101 && y_pointer == 23)
||(x_pointer == 102 && y_pointer == 23)
||(x_pointer == 103 && y_pointer == 23)
||(x_pointer == 104 && y_pointer == 23)
||(x_pointer == 105 && y_pointer == 23)
||(x_pointer == 106 && y_pointer == 23)
||(x_pointer == 107 && y_pointer == 23)
||(x_pointer == 108 && y_pointer == 23)
||(x_pointer == 109 && y_pointer == 23)
||(x_pointer == 110 && y_pointer == 23)
||(x_pointer == 111 && y_pointer == 23)
||(x_pointer == 112 && y_pointer == 23)
||(x_pointer == 155 && y_pointer == 23)
||(x_pointer == 156 && y_pointer == 23)
||(x_pointer == 157 && y_pointer == 23)
||(x_pointer == 2 && y_pointer == 24)
||(x_pointer == 3 && y_pointer == 24)
||(x_pointer == 4 && y_pointer == 24)
||(x_pointer == 50 && y_pointer == 24)
||(x_pointer == 51 && y_pointer == 24)
||(x_pointer == 52 && y_pointer == 24)
||(x_pointer == 53 && y_pointer == 24)
||(x_pointer == 54 && y_pointer == 24)
||(x_pointer == 55 && y_pointer == 24)
||(x_pointer == 56 && y_pointer == 24)
||(x_pointer == 57 && y_pointer == 24)
||(x_pointer == 58 && y_pointer == 24)
||(x_pointer == 59 && y_pointer == 24)
||(x_pointer == 60 && y_pointer == 24)
||(x_pointer == 61 && y_pointer == 24)
||(x_pointer == 62 && y_pointer == 24)
||(x_pointer == 63 && y_pointer == 24)
||(x_pointer == 64 && y_pointer == 24)
||(x_pointer == 65 && y_pointer == 24)
||(x_pointer == 66 && y_pointer == 24)
||(x_pointer == 67 && y_pointer == 24)
||(x_pointer == 68 && y_pointer == 24)
||(x_pointer == 69 && y_pointer == 24)
||(x_pointer == 70 && y_pointer == 24)
||(x_pointer == 71 && y_pointer == 24)
||(x_pointer == 72 && y_pointer == 24)
||(x_pointer == 73 && y_pointer == 24)
||(x_pointer == 89 && y_pointer == 24)
||(x_pointer == 90 && y_pointer == 24)
||(x_pointer == 91 && y_pointer == 24)
||(x_pointer == 92 && y_pointer == 24)
||(x_pointer == 93 && y_pointer == 24)
||(x_pointer == 94 && y_pointer == 24)
||(x_pointer == 95 && y_pointer == 24)
||(x_pointer == 96 && y_pointer == 24)
||(x_pointer == 97 && y_pointer == 24)
||(x_pointer == 98 && y_pointer == 24)
||(x_pointer == 99 && y_pointer == 24)
||(x_pointer == 100 && y_pointer == 24)
||(x_pointer == 101 && y_pointer == 24)
||(x_pointer == 102 && y_pointer == 24)
||(x_pointer == 103 && y_pointer == 24)
||(x_pointer == 104 && y_pointer == 24)
||(x_pointer == 105 && y_pointer == 24)
||(x_pointer == 106 && y_pointer == 24)
||(x_pointer == 107 && y_pointer == 24)
||(x_pointer == 108 && y_pointer == 24)
||(x_pointer == 109 && y_pointer == 24)
||(x_pointer == 110 && y_pointer == 24)
||(x_pointer == 111 && y_pointer == 24)
||(x_pointer == 112 && y_pointer == 24)
||(x_pointer == 155 && y_pointer == 24)
||(x_pointer == 156 && y_pointer == 24)
||(x_pointer == 157 && y_pointer == 24)
||(x_pointer == 2 && y_pointer == 25)
||(x_pointer == 3 && y_pointer == 25)
||(x_pointer == 4 && y_pointer == 25)
||(x_pointer == 50 && y_pointer == 25)
||(x_pointer == 51 && y_pointer == 25)
||(x_pointer == 52 && y_pointer == 25)
||(x_pointer == 53 && y_pointer == 25)
||(x_pointer == 54 && y_pointer == 25)
||(x_pointer == 55 && y_pointer == 25)
||(x_pointer == 56 && y_pointer == 25)
||(x_pointer == 57 && y_pointer == 25)
||(x_pointer == 58 && y_pointer == 25)
||(x_pointer == 59 && y_pointer == 25)
||(x_pointer == 60 && y_pointer == 25)
||(x_pointer == 61 && y_pointer == 25)
||(x_pointer == 62 && y_pointer == 25)
||(x_pointer == 63 && y_pointer == 25)
||(x_pointer == 64 && y_pointer == 25)
||(x_pointer == 65 && y_pointer == 25)
||(x_pointer == 66 && y_pointer == 25)
||(x_pointer == 67 && y_pointer == 25)
||(x_pointer == 68 && y_pointer == 25)
||(x_pointer == 69 && y_pointer == 25)
||(x_pointer == 70 && y_pointer == 25)
||(x_pointer == 71 && y_pointer == 25)
||(x_pointer == 72 && y_pointer == 25)
||(x_pointer == 73 && y_pointer == 25)
||(x_pointer == 89 && y_pointer == 25)
||(x_pointer == 90 && y_pointer == 25)
||(x_pointer == 91 && y_pointer == 25)
||(x_pointer == 92 && y_pointer == 25)
||(x_pointer == 93 && y_pointer == 25)
||(x_pointer == 94 && y_pointer == 25)
||(x_pointer == 95 && y_pointer == 25)
||(x_pointer == 96 && y_pointer == 25)
||(x_pointer == 97 && y_pointer == 25)
||(x_pointer == 98 && y_pointer == 25)
||(x_pointer == 99 && y_pointer == 25)
||(x_pointer == 100 && y_pointer == 25)
||(x_pointer == 101 && y_pointer == 25)
||(x_pointer == 102 && y_pointer == 25)
||(x_pointer == 103 && y_pointer == 25)
||(x_pointer == 104 && y_pointer == 25)
||(x_pointer == 105 && y_pointer == 25)
||(x_pointer == 106 && y_pointer == 25)
||(x_pointer == 107 && y_pointer == 25)
||(x_pointer == 108 && y_pointer == 25)
||(x_pointer == 109 && y_pointer == 25)
||(x_pointer == 110 && y_pointer == 25)
||(x_pointer == 111 && y_pointer == 25)
||(x_pointer == 112 && y_pointer == 25)
||(x_pointer == 155 && y_pointer == 25)
||(x_pointer == 156 && y_pointer == 25)
||(x_pointer == 157 && y_pointer == 25)
||(x_pointer == 2 && y_pointer == 26)
||(x_pointer == 3 && y_pointer == 26)
||(x_pointer == 4 && y_pointer == 26)
||(x_pointer == 50 && y_pointer == 26)
||(x_pointer == 51 && y_pointer == 26)
||(x_pointer == 52 && y_pointer == 26)
||(x_pointer == 53 && y_pointer == 26)
||(x_pointer == 54 && y_pointer == 26)
||(x_pointer == 55 && y_pointer == 26)
||(x_pointer == 56 && y_pointer == 26)
||(x_pointer == 57 && y_pointer == 26)
||(x_pointer == 58 && y_pointer == 26)
||(x_pointer == 59 && y_pointer == 26)
||(x_pointer == 60 && y_pointer == 26)
||(x_pointer == 61 && y_pointer == 26)
||(x_pointer == 62 && y_pointer == 26)
||(x_pointer == 63 && y_pointer == 26)
||(x_pointer == 64 && y_pointer == 26)
||(x_pointer == 65 && y_pointer == 26)
||(x_pointer == 66 && y_pointer == 26)
||(x_pointer == 67 && y_pointer == 26)
||(x_pointer == 68 && y_pointer == 26)
||(x_pointer == 69 && y_pointer == 26)
||(x_pointer == 70 && y_pointer == 26)
||(x_pointer == 71 && y_pointer == 26)
||(x_pointer == 72 && y_pointer == 26)
||(x_pointer == 73 && y_pointer == 26)
||(x_pointer == 89 && y_pointer == 26)
||(x_pointer == 90 && y_pointer == 26)
||(x_pointer == 91 && y_pointer == 26)
||(x_pointer == 92 && y_pointer == 26)
||(x_pointer == 93 && y_pointer == 26)
||(x_pointer == 94 && y_pointer == 26)
||(x_pointer == 95 && y_pointer == 26)
||(x_pointer == 96 && y_pointer == 26)
||(x_pointer == 97 && y_pointer == 26)
||(x_pointer == 98 && y_pointer == 26)
||(x_pointer == 99 && y_pointer == 26)
||(x_pointer == 100 && y_pointer == 26)
||(x_pointer == 101 && y_pointer == 26)
||(x_pointer == 102 && y_pointer == 26)
||(x_pointer == 103 && y_pointer == 26)
||(x_pointer == 104 && y_pointer == 26)
||(x_pointer == 105 && y_pointer == 26)
||(x_pointer == 106 && y_pointer == 26)
||(x_pointer == 107 && y_pointer == 26)
||(x_pointer == 108 && y_pointer == 26)
||(x_pointer == 109 && y_pointer == 26)
||(x_pointer == 110 && y_pointer == 26)
||(x_pointer == 111 && y_pointer == 26)
||(x_pointer == 112 && y_pointer == 26)
||(x_pointer == 155 && y_pointer == 26)
||(x_pointer == 156 && y_pointer == 26)
||(x_pointer == 157 && y_pointer == 26)
||(x_pointer == 2 && y_pointer == 27)
||(x_pointer == 3 && y_pointer == 27)
||(x_pointer == 4 && y_pointer == 27)
||(x_pointer == 50 && y_pointer == 27)
||(x_pointer == 51 && y_pointer == 27)
||(x_pointer == 52 && y_pointer == 27)
||(x_pointer == 53 && y_pointer == 27)
||(x_pointer == 54 && y_pointer == 27)
||(x_pointer == 55 && y_pointer == 27)
||(x_pointer == 56 && y_pointer == 27)
||(x_pointer == 57 && y_pointer == 27)
||(x_pointer == 58 && y_pointer == 27)
||(x_pointer == 59 && y_pointer == 27)
||(x_pointer == 60 && y_pointer == 27)
||(x_pointer == 61 && y_pointer == 27)
||(x_pointer == 62 && y_pointer == 27)
||(x_pointer == 63 && y_pointer == 27)
||(x_pointer == 64 && y_pointer == 27)
||(x_pointer == 65 && y_pointer == 27)
||(x_pointer == 66 && y_pointer == 27)
||(x_pointer == 67 && y_pointer == 27)
||(x_pointer == 68 && y_pointer == 27)
||(x_pointer == 69 && y_pointer == 27)
||(x_pointer == 70 && y_pointer == 27)
||(x_pointer == 71 && y_pointer == 27)
||(x_pointer == 72 && y_pointer == 27)
||(x_pointer == 73 && y_pointer == 27)
||(x_pointer == 89 && y_pointer == 27)
||(x_pointer == 90 && y_pointer == 27)
||(x_pointer == 91 && y_pointer == 27)
||(x_pointer == 92 && y_pointer == 27)
||(x_pointer == 93 && y_pointer == 27)
||(x_pointer == 94 && y_pointer == 27)
||(x_pointer == 95 && y_pointer == 27)
||(x_pointer == 96 && y_pointer == 27)
||(x_pointer == 97 && y_pointer == 27)
||(x_pointer == 98 && y_pointer == 27)
||(x_pointer == 99 && y_pointer == 27)
||(x_pointer == 100 && y_pointer == 27)
||(x_pointer == 101 && y_pointer == 27)
||(x_pointer == 102 && y_pointer == 27)
||(x_pointer == 103 && y_pointer == 27)
||(x_pointer == 104 && y_pointer == 27)
||(x_pointer == 105 && y_pointer == 27)
||(x_pointer == 106 && y_pointer == 27)
||(x_pointer == 107 && y_pointer == 27)
||(x_pointer == 108 && y_pointer == 27)
||(x_pointer == 109 && y_pointer == 27)
||(x_pointer == 110 && y_pointer == 27)
||(x_pointer == 111 && y_pointer == 27)
||(x_pointer == 112 && y_pointer == 27)
||(x_pointer == 155 && y_pointer == 27)
||(x_pointer == 156 && y_pointer == 27)
||(x_pointer == 157 && y_pointer == 27)
||(x_pointer == 2 && y_pointer == 28)
||(x_pointer == 3 && y_pointer == 28)
||(x_pointer == 4 && y_pointer == 28)
||(x_pointer == 50 && y_pointer == 28)
||(x_pointer == 51 && y_pointer == 28)
||(x_pointer == 52 && y_pointer == 28)
||(x_pointer == 53 && y_pointer == 28)
||(x_pointer == 54 && y_pointer == 28)
||(x_pointer == 55 && y_pointer == 28)
||(x_pointer == 56 && y_pointer == 28)
||(x_pointer == 57 && y_pointer == 28)
||(x_pointer == 58 && y_pointer == 28)
||(x_pointer == 59 && y_pointer == 28)
||(x_pointer == 60 && y_pointer == 28)
||(x_pointer == 61 && y_pointer == 28)
||(x_pointer == 62 && y_pointer == 28)
||(x_pointer == 63 && y_pointer == 28)
||(x_pointer == 64 && y_pointer == 28)
||(x_pointer == 65 && y_pointer == 28)
||(x_pointer == 66 && y_pointer == 28)
||(x_pointer == 67 && y_pointer == 28)
||(x_pointer == 68 && y_pointer == 28)
||(x_pointer == 69 && y_pointer == 28)
||(x_pointer == 70 && y_pointer == 28)
||(x_pointer == 71 && y_pointer == 28)
||(x_pointer == 72 && y_pointer == 28)
||(x_pointer == 73 && y_pointer == 28)
||(x_pointer == 89 && y_pointer == 28)
||(x_pointer == 90 && y_pointer == 28)
||(x_pointer == 91 && y_pointer == 28)
||(x_pointer == 92 && y_pointer == 28)
||(x_pointer == 93 && y_pointer == 28)
||(x_pointer == 94 && y_pointer == 28)
||(x_pointer == 95 && y_pointer == 28)
||(x_pointer == 96 && y_pointer == 28)
||(x_pointer == 97 && y_pointer == 28)
||(x_pointer == 98 && y_pointer == 28)
||(x_pointer == 99 && y_pointer == 28)
||(x_pointer == 100 && y_pointer == 28)
||(x_pointer == 101 && y_pointer == 28)
||(x_pointer == 102 && y_pointer == 28)
||(x_pointer == 103 && y_pointer == 28)
||(x_pointer == 104 && y_pointer == 28)
||(x_pointer == 105 && y_pointer == 28)
||(x_pointer == 106 && y_pointer == 28)
||(x_pointer == 107 && y_pointer == 28)
||(x_pointer == 108 && y_pointer == 28)
||(x_pointer == 109 && y_pointer == 28)
||(x_pointer == 110 && y_pointer == 28)
||(x_pointer == 111 && y_pointer == 28)
||(x_pointer == 112 && y_pointer == 28)
||(x_pointer == 155 && y_pointer == 28)
||(x_pointer == 156 && y_pointer == 28)
||(x_pointer == 157 && y_pointer == 28)
||(x_pointer == 2 && y_pointer == 29)
||(x_pointer == 3 && y_pointer == 29)
||(x_pointer == 4 && y_pointer == 29)
||(x_pointer == 50 && y_pointer == 29)
||(x_pointer == 51 && y_pointer == 29)
||(x_pointer == 52 && y_pointer == 29)
||(x_pointer == 53 && y_pointer == 29)
||(x_pointer == 54 && y_pointer == 29)
||(x_pointer == 55 && y_pointer == 29)
||(x_pointer == 56 && y_pointer == 29)
||(x_pointer == 57 && y_pointer == 29)
||(x_pointer == 58 && y_pointer == 29)
||(x_pointer == 59 && y_pointer == 29)
||(x_pointer == 60 && y_pointer == 29)
||(x_pointer == 61 && y_pointer == 29)
||(x_pointer == 62 && y_pointer == 29)
||(x_pointer == 63 && y_pointer == 29)
||(x_pointer == 64 && y_pointer == 29)
||(x_pointer == 65 && y_pointer == 29)
||(x_pointer == 66 && y_pointer == 29)
||(x_pointer == 67 && y_pointer == 29)
||(x_pointer == 68 && y_pointer == 29)
||(x_pointer == 69 && y_pointer == 29)
||(x_pointer == 70 && y_pointer == 29)
||(x_pointer == 71 && y_pointer == 29)
||(x_pointer == 72 && y_pointer == 29)
||(x_pointer == 73 && y_pointer == 29)
||(x_pointer == 89 && y_pointer == 29)
||(x_pointer == 90 && y_pointer == 29)
||(x_pointer == 91 && y_pointer == 29)
||(x_pointer == 92 && y_pointer == 29)
||(x_pointer == 93 && y_pointer == 29)
||(x_pointer == 94 && y_pointer == 29)
||(x_pointer == 95 && y_pointer == 29)
||(x_pointer == 96 && y_pointer == 29)
||(x_pointer == 97 && y_pointer == 29)
||(x_pointer == 98 && y_pointer == 29)
||(x_pointer == 99 && y_pointer == 29)
||(x_pointer == 100 && y_pointer == 29)
||(x_pointer == 101 && y_pointer == 29)
||(x_pointer == 102 && y_pointer == 29)
||(x_pointer == 103 && y_pointer == 29)
||(x_pointer == 104 && y_pointer == 29)
||(x_pointer == 105 && y_pointer == 29)
||(x_pointer == 106 && y_pointer == 29)
||(x_pointer == 107 && y_pointer == 29)
||(x_pointer == 108 && y_pointer == 29)
||(x_pointer == 109 && y_pointer == 29)
||(x_pointer == 110 && y_pointer == 29)
||(x_pointer == 111 && y_pointer == 29)
||(x_pointer == 112 && y_pointer == 29)
||(x_pointer == 155 && y_pointer == 29)
||(x_pointer == 156 && y_pointer == 29)
||(x_pointer == 157 && y_pointer == 29)
||(x_pointer == 2 && y_pointer == 30)
||(x_pointer == 3 && y_pointer == 30)
||(x_pointer == 4 && y_pointer == 30)
||(x_pointer == 50 && y_pointer == 30)
||(x_pointer == 51 && y_pointer == 30)
||(x_pointer == 52 && y_pointer == 30)
||(x_pointer == 53 && y_pointer == 30)
||(x_pointer == 54 && y_pointer == 30)
||(x_pointer == 55 && y_pointer == 30)
||(x_pointer == 56 && y_pointer == 30)
||(x_pointer == 57 && y_pointer == 30)
||(x_pointer == 58 && y_pointer == 30)
||(x_pointer == 59 && y_pointer == 30)
||(x_pointer == 60 && y_pointer == 30)
||(x_pointer == 61 && y_pointer == 30)
||(x_pointer == 62 && y_pointer == 30)
||(x_pointer == 63 && y_pointer == 30)
||(x_pointer == 64 && y_pointer == 30)
||(x_pointer == 65 && y_pointer == 30)
||(x_pointer == 66 && y_pointer == 30)
||(x_pointer == 67 && y_pointer == 30)
||(x_pointer == 68 && y_pointer == 30)
||(x_pointer == 69 && y_pointer == 30)
||(x_pointer == 70 && y_pointer == 30)
||(x_pointer == 71 && y_pointer == 30)
||(x_pointer == 72 && y_pointer == 30)
||(x_pointer == 73 && y_pointer == 30)
||(x_pointer == 89 && y_pointer == 30)
||(x_pointer == 90 && y_pointer == 30)
||(x_pointer == 91 && y_pointer == 30)
||(x_pointer == 92 && y_pointer == 30)
||(x_pointer == 93 && y_pointer == 30)
||(x_pointer == 94 && y_pointer == 30)
||(x_pointer == 95 && y_pointer == 30)
||(x_pointer == 96 && y_pointer == 30)
||(x_pointer == 97 && y_pointer == 30)
||(x_pointer == 98 && y_pointer == 30)
||(x_pointer == 99 && y_pointer == 30)
||(x_pointer == 100 && y_pointer == 30)
||(x_pointer == 101 && y_pointer == 30)
||(x_pointer == 102 && y_pointer == 30)
||(x_pointer == 103 && y_pointer == 30)
||(x_pointer == 104 && y_pointer == 30)
||(x_pointer == 105 && y_pointer == 30)
||(x_pointer == 106 && y_pointer == 30)
||(x_pointer == 107 && y_pointer == 30)
||(x_pointer == 108 && y_pointer == 30)
||(x_pointer == 109 && y_pointer == 30)
||(x_pointer == 110 && y_pointer == 30)
||(x_pointer == 111 && y_pointer == 30)
||(x_pointer == 112 && y_pointer == 30)
||(x_pointer == 155 && y_pointer == 30)
||(x_pointer == 156 && y_pointer == 30)
||(x_pointer == 157 && y_pointer == 30)
||(x_pointer == 2 && y_pointer == 31)
||(x_pointer == 3 && y_pointer == 31)
||(x_pointer == 4 && y_pointer == 31)
||(x_pointer == 50 && y_pointer == 31)
||(x_pointer == 51 && y_pointer == 31)
||(x_pointer == 52 && y_pointer == 31)
||(x_pointer == 53 && y_pointer == 31)
||(x_pointer == 54 && y_pointer == 31)
||(x_pointer == 55 && y_pointer == 31)
||(x_pointer == 56 && y_pointer == 31)
||(x_pointer == 57 && y_pointer == 31)
||(x_pointer == 58 && y_pointer == 31)
||(x_pointer == 59 && y_pointer == 31)
||(x_pointer == 60 && y_pointer == 31)
||(x_pointer == 61 && y_pointer == 31)
||(x_pointer == 62 && y_pointer == 31)
||(x_pointer == 63 && y_pointer == 31)
||(x_pointer == 64 && y_pointer == 31)
||(x_pointer == 65 && y_pointer == 31)
||(x_pointer == 66 && y_pointer == 31)
||(x_pointer == 67 && y_pointer == 31)
||(x_pointer == 68 && y_pointer == 31)
||(x_pointer == 69 && y_pointer == 31)
||(x_pointer == 70 && y_pointer == 31)
||(x_pointer == 71 && y_pointer == 31)
||(x_pointer == 72 && y_pointer == 31)
||(x_pointer == 73 && y_pointer == 31)
||(x_pointer == 89 && y_pointer == 31)
||(x_pointer == 90 && y_pointer == 31)
||(x_pointer == 91 && y_pointer == 31)
||(x_pointer == 92 && y_pointer == 31)
||(x_pointer == 93 && y_pointer == 31)
||(x_pointer == 94 && y_pointer == 31)
||(x_pointer == 95 && y_pointer == 31)
||(x_pointer == 96 && y_pointer == 31)
||(x_pointer == 97 && y_pointer == 31)
||(x_pointer == 98 && y_pointer == 31)
||(x_pointer == 99 && y_pointer == 31)
||(x_pointer == 100 && y_pointer == 31)
||(x_pointer == 101 && y_pointer == 31)
||(x_pointer == 102 && y_pointer == 31)
||(x_pointer == 103 && y_pointer == 31)
||(x_pointer == 104 && y_pointer == 31)
||(x_pointer == 105 && y_pointer == 31)
||(x_pointer == 106 && y_pointer == 31)
||(x_pointer == 107 && y_pointer == 31)
||(x_pointer == 108 && y_pointer == 31)
||(x_pointer == 109 && y_pointer == 31)
||(x_pointer == 110 && y_pointer == 31)
||(x_pointer == 111 && y_pointer == 31)
||(x_pointer == 112 && y_pointer == 31)
||(x_pointer == 155 && y_pointer == 31)
||(x_pointer == 156 && y_pointer == 31)
||(x_pointer == 157 && y_pointer == 31)
||(x_pointer == 2 && y_pointer == 32)
||(x_pointer == 3 && y_pointer == 32)
||(x_pointer == 4 && y_pointer == 32)
||(x_pointer == 50 && y_pointer == 32)
||(x_pointer == 51 && y_pointer == 32)
||(x_pointer == 52 && y_pointer == 32)
||(x_pointer == 53 && y_pointer == 32)
||(x_pointer == 54 && y_pointer == 32)
||(x_pointer == 55 && y_pointer == 32)
||(x_pointer == 56 && y_pointer == 32)
||(x_pointer == 57 && y_pointer == 32)
||(x_pointer == 58 && y_pointer == 32)
||(x_pointer == 59 && y_pointer == 32)
||(x_pointer == 60 && y_pointer == 32)
||(x_pointer == 61 && y_pointer == 32)
||(x_pointer == 62 && y_pointer == 32)
||(x_pointer == 63 && y_pointer == 32)
||(x_pointer == 64 && y_pointer == 32)
||(x_pointer == 65 && y_pointer == 32)
||(x_pointer == 66 && y_pointer == 32)
||(x_pointer == 67 && y_pointer == 32)
||(x_pointer == 68 && y_pointer == 32)
||(x_pointer == 69 && y_pointer == 32)
||(x_pointer == 70 && y_pointer == 32)
||(x_pointer == 71 && y_pointer == 32)
||(x_pointer == 72 && y_pointer == 32)
||(x_pointer == 73 && y_pointer == 32)
||(x_pointer == 89 && y_pointer == 32)
||(x_pointer == 90 && y_pointer == 32)
||(x_pointer == 91 && y_pointer == 32)
||(x_pointer == 92 && y_pointer == 32)
||(x_pointer == 93 && y_pointer == 32)
||(x_pointer == 94 && y_pointer == 32)
||(x_pointer == 95 && y_pointer == 32)
||(x_pointer == 96 && y_pointer == 32)
||(x_pointer == 97 && y_pointer == 32)
||(x_pointer == 98 && y_pointer == 32)
||(x_pointer == 99 && y_pointer == 32)
||(x_pointer == 100 && y_pointer == 32)
||(x_pointer == 101 && y_pointer == 32)
||(x_pointer == 102 && y_pointer == 32)
||(x_pointer == 103 && y_pointer == 32)
||(x_pointer == 104 && y_pointer == 32)
||(x_pointer == 105 && y_pointer == 32)
||(x_pointer == 106 && y_pointer == 32)
||(x_pointer == 107 && y_pointer == 32)
||(x_pointer == 108 && y_pointer == 32)
||(x_pointer == 109 && y_pointer == 32)
||(x_pointer == 110 && y_pointer == 32)
||(x_pointer == 111 && y_pointer == 32)
||(x_pointer == 112 && y_pointer == 32)
||(x_pointer == 155 && y_pointer == 32)
||(x_pointer == 156 && y_pointer == 32)
||(x_pointer == 157 && y_pointer == 32)
||(x_pointer == 2 && y_pointer == 33)
||(x_pointer == 3 && y_pointer == 33)
||(x_pointer == 4 && y_pointer == 33)
||(x_pointer == 50 && y_pointer == 33)
||(x_pointer == 51 && y_pointer == 33)
||(x_pointer == 52 && y_pointer == 33)
||(x_pointer == 53 && y_pointer == 33)
||(x_pointer == 54 && y_pointer == 33)
||(x_pointer == 55 && y_pointer == 33)
||(x_pointer == 56 && y_pointer == 33)
||(x_pointer == 57 && y_pointer == 33)
||(x_pointer == 58 && y_pointer == 33)
||(x_pointer == 59 && y_pointer == 33)
||(x_pointer == 60 && y_pointer == 33)
||(x_pointer == 61 && y_pointer == 33)
||(x_pointer == 62 && y_pointer == 33)
||(x_pointer == 63 && y_pointer == 33)
||(x_pointer == 64 && y_pointer == 33)
||(x_pointer == 65 && y_pointer == 33)
||(x_pointer == 66 && y_pointer == 33)
||(x_pointer == 67 && y_pointer == 33)
||(x_pointer == 68 && y_pointer == 33)
||(x_pointer == 69 && y_pointer == 33)
||(x_pointer == 70 && y_pointer == 33)
||(x_pointer == 71 && y_pointer == 33)
||(x_pointer == 72 && y_pointer == 33)
||(x_pointer == 73 && y_pointer == 33)
||(x_pointer == 89 && y_pointer == 33)
||(x_pointer == 90 && y_pointer == 33)
||(x_pointer == 91 && y_pointer == 33)
||(x_pointer == 92 && y_pointer == 33)
||(x_pointer == 93 && y_pointer == 33)
||(x_pointer == 94 && y_pointer == 33)
||(x_pointer == 95 && y_pointer == 33)
||(x_pointer == 96 && y_pointer == 33)
||(x_pointer == 97 && y_pointer == 33)
||(x_pointer == 98 && y_pointer == 33)
||(x_pointer == 99 && y_pointer == 33)
||(x_pointer == 100 && y_pointer == 33)
||(x_pointer == 101 && y_pointer == 33)
||(x_pointer == 102 && y_pointer == 33)
||(x_pointer == 103 && y_pointer == 33)
||(x_pointer == 104 && y_pointer == 33)
||(x_pointer == 105 && y_pointer == 33)
||(x_pointer == 106 && y_pointer == 33)
||(x_pointer == 107 && y_pointer == 33)
||(x_pointer == 108 && y_pointer == 33)
||(x_pointer == 109 && y_pointer == 33)
||(x_pointer == 110 && y_pointer == 33)
||(x_pointer == 111 && y_pointer == 33)
||(x_pointer == 112 && y_pointer == 33)
||(x_pointer == 155 && y_pointer == 33)
||(x_pointer == 156 && y_pointer == 33)
||(x_pointer == 157 && y_pointer == 33)
||(x_pointer == 2 && y_pointer == 34)
||(x_pointer == 3 && y_pointer == 34)
||(x_pointer == 4 && y_pointer == 34)
||(x_pointer == 50 && y_pointer == 34)
||(x_pointer == 51 && y_pointer == 34)
||(x_pointer == 52 && y_pointer == 34)
||(x_pointer == 53 && y_pointer == 34)
||(x_pointer == 54 && y_pointer == 34)
||(x_pointer == 55 && y_pointer == 34)
||(x_pointer == 56 && y_pointer == 34)
||(x_pointer == 57 && y_pointer == 34)
||(x_pointer == 58 && y_pointer == 34)
||(x_pointer == 59 && y_pointer == 34)
||(x_pointer == 60 && y_pointer == 34)
||(x_pointer == 61 && y_pointer == 34)
||(x_pointer == 62 && y_pointer == 34)
||(x_pointer == 63 && y_pointer == 34)
||(x_pointer == 64 && y_pointer == 34)
||(x_pointer == 65 && y_pointer == 34)
||(x_pointer == 66 && y_pointer == 34)
||(x_pointer == 67 && y_pointer == 34)
||(x_pointer == 68 && y_pointer == 34)
||(x_pointer == 69 && y_pointer == 34)
||(x_pointer == 70 && y_pointer == 34)
||(x_pointer == 71 && y_pointer == 34)
||(x_pointer == 72 && y_pointer == 34)
||(x_pointer == 73 && y_pointer == 34)
||(x_pointer == 89 && y_pointer == 34)
||(x_pointer == 90 && y_pointer == 34)
||(x_pointer == 91 && y_pointer == 34)
||(x_pointer == 92 && y_pointer == 34)
||(x_pointer == 93 && y_pointer == 34)
||(x_pointer == 94 && y_pointer == 34)
||(x_pointer == 95 && y_pointer == 34)
||(x_pointer == 96 && y_pointer == 34)
||(x_pointer == 97 && y_pointer == 34)
||(x_pointer == 98 && y_pointer == 34)
||(x_pointer == 99 && y_pointer == 34)
||(x_pointer == 100 && y_pointer == 34)
||(x_pointer == 101 && y_pointer == 34)
||(x_pointer == 102 && y_pointer == 34)
||(x_pointer == 103 && y_pointer == 34)
||(x_pointer == 104 && y_pointer == 34)
||(x_pointer == 105 && y_pointer == 34)
||(x_pointer == 106 && y_pointer == 34)
||(x_pointer == 107 && y_pointer == 34)
||(x_pointer == 108 && y_pointer == 34)
||(x_pointer == 109 && y_pointer == 34)
||(x_pointer == 110 && y_pointer == 34)
||(x_pointer == 111 && y_pointer == 34)
||(x_pointer == 112 && y_pointer == 34)
||(x_pointer == 155 && y_pointer == 34)
||(x_pointer == 156 && y_pointer == 34)
||(x_pointer == 157 && y_pointer == 34)
||(x_pointer == 2 && y_pointer == 35)
||(x_pointer == 3 && y_pointer == 35)
||(x_pointer == 4 && y_pointer == 35)
||(x_pointer == 50 && y_pointer == 35)
||(x_pointer == 51 && y_pointer == 35)
||(x_pointer == 52 && y_pointer == 35)
||(x_pointer == 53 && y_pointer == 35)
||(x_pointer == 54 && y_pointer == 35)
||(x_pointer == 55 && y_pointer == 35)
||(x_pointer == 56 && y_pointer == 35)
||(x_pointer == 57 && y_pointer == 35)
||(x_pointer == 58 && y_pointer == 35)
||(x_pointer == 59 && y_pointer == 35)
||(x_pointer == 60 && y_pointer == 35)
||(x_pointer == 61 && y_pointer == 35)
||(x_pointer == 62 && y_pointer == 35)
||(x_pointer == 63 && y_pointer == 35)
||(x_pointer == 64 && y_pointer == 35)
||(x_pointer == 65 && y_pointer == 35)
||(x_pointer == 66 && y_pointer == 35)
||(x_pointer == 67 && y_pointer == 35)
||(x_pointer == 68 && y_pointer == 35)
||(x_pointer == 69 && y_pointer == 35)
||(x_pointer == 70 && y_pointer == 35)
||(x_pointer == 71 && y_pointer == 35)
||(x_pointer == 72 && y_pointer == 35)
||(x_pointer == 73 && y_pointer == 35)
||(x_pointer == 89 && y_pointer == 35)
||(x_pointer == 90 && y_pointer == 35)
||(x_pointer == 91 && y_pointer == 35)
||(x_pointer == 92 && y_pointer == 35)
||(x_pointer == 93 && y_pointer == 35)
||(x_pointer == 94 && y_pointer == 35)
||(x_pointer == 95 && y_pointer == 35)
||(x_pointer == 96 && y_pointer == 35)
||(x_pointer == 97 && y_pointer == 35)
||(x_pointer == 98 && y_pointer == 35)
||(x_pointer == 99 && y_pointer == 35)
||(x_pointer == 100 && y_pointer == 35)
||(x_pointer == 101 && y_pointer == 35)
||(x_pointer == 102 && y_pointer == 35)
||(x_pointer == 103 && y_pointer == 35)
||(x_pointer == 104 && y_pointer == 35)
||(x_pointer == 105 && y_pointer == 35)
||(x_pointer == 106 && y_pointer == 35)
||(x_pointer == 107 && y_pointer == 35)
||(x_pointer == 108 && y_pointer == 35)
||(x_pointer == 109 && y_pointer == 35)
||(x_pointer == 110 && y_pointer == 35)
||(x_pointer == 111 && y_pointer == 35)
||(x_pointer == 112 && y_pointer == 35)
||(x_pointer == 155 && y_pointer == 35)
||(x_pointer == 156 && y_pointer == 35)
||(x_pointer == 157 && y_pointer == 35)
||(x_pointer == 2 && y_pointer == 36)
||(x_pointer == 3 && y_pointer == 36)
||(x_pointer == 4 && y_pointer == 36)
||(x_pointer == 50 && y_pointer == 36)
||(x_pointer == 51 && y_pointer == 36)
||(x_pointer == 52 && y_pointer == 36)
||(x_pointer == 53 && y_pointer == 36)
||(x_pointer == 54 && y_pointer == 36)
||(x_pointer == 55 && y_pointer == 36)
||(x_pointer == 56 && y_pointer == 36)
||(x_pointer == 57 && y_pointer == 36)
||(x_pointer == 58 && y_pointer == 36)
||(x_pointer == 59 && y_pointer == 36)
||(x_pointer == 60 && y_pointer == 36)
||(x_pointer == 61 && y_pointer == 36)
||(x_pointer == 62 && y_pointer == 36)
||(x_pointer == 63 && y_pointer == 36)
||(x_pointer == 64 && y_pointer == 36)
||(x_pointer == 65 && y_pointer == 36)
||(x_pointer == 66 && y_pointer == 36)
||(x_pointer == 67 && y_pointer == 36)
||(x_pointer == 68 && y_pointer == 36)
||(x_pointer == 69 && y_pointer == 36)
||(x_pointer == 70 && y_pointer == 36)
||(x_pointer == 71 && y_pointer == 36)
||(x_pointer == 72 && y_pointer == 36)
||(x_pointer == 73 && y_pointer == 36)
||(x_pointer == 89 && y_pointer == 36)
||(x_pointer == 90 && y_pointer == 36)
||(x_pointer == 91 && y_pointer == 36)
||(x_pointer == 92 && y_pointer == 36)
||(x_pointer == 93 && y_pointer == 36)
||(x_pointer == 94 && y_pointer == 36)
||(x_pointer == 95 && y_pointer == 36)
||(x_pointer == 96 && y_pointer == 36)
||(x_pointer == 97 && y_pointer == 36)
||(x_pointer == 98 && y_pointer == 36)
||(x_pointer == 99 && y_pointer == 36)
||(x_pointer == 100 && y_pointer == 36)
||(x_pointer == 101 && y_pointer == 36)
||(x_pointer == 102 && y_pointer == 36)
||(x_pointer == 103 && y_pointer == 36)
||(x_pointer == 104 && y_pointer == 36)
||(x_pointer == 105 && y_pointer == 36)
||(x_pointer == 106 && y_pointer == 36)
||(x_pointer == 107 && y_pointer == 36)
||(x_pointer == 108 && y_pointer == 36)
||(x_pointer == 109 && y_pointer == 36)
||(x_pointer == 110 && y_pointer == 36)
||(x_pointer == 111 && y_pointer == 36)
||(x_pointer == 112 && y_pointer == 36)
||(x_pointer == 155 && y_pointer == 36)
||(x_pointer == 156 && y_pointer == 36)
||(x_pointer == 157 && y_pointer == 36)
||(x_pointer == 2 && y_pointer == 37)
||(x_pointer == 3 && y_pointer == 37)
||(x_pointer == 4 && y_pointer == 37)
||(x_pointer == 50 && y_pointer == 37)
||(x_pointer == 51 && y_pointer == 37)
||(x_pointer == 52 && y_pointer == 37)
||(x_pointer == 53 && y_pointer == 37)
||(x_pointer == 54 && y_pointer == 37)
||(x_pointer == 55 && y_pointer == 37)
||(x_pointer == 56 && y_pointer == 37)
||(x_pointer == 57 && y_pointer == 37)
||(x_pointer == 58 && y_pointer == 37)
||(x_pointer == 59 && y_pointer == 37)
||(x_pointer == 60 && y_pointer == 37)
||(x_pointer == 61 && y_pointer == 37)
||(x_pointer == 62 && y_pointer == 37)
||(x_pointer == 63 && y_pointer == 37)
||(x_pointer == 64 && y_pointer == 37)
||(x_pointer == 65 && y_pointer == 37)
||(x_pointer == 66 && y_pointer == 37)
||(x_pointer == 67 && y_pointer == 37)
||(x_pointer == 68 && y_pointer == 37)
||(x_pointer == 69 && y_pointer == 37)
||(x_pointer == 70 && y_pointer == 37)
||(x_pointer == 71 && y_pointer == 37)
||(x_pointer == 72 && y_pointer == 37)
||(x_pointer == 73 && y_pointer == 37)
||(x_pointer == 89 && y_pointer == 37)
||(x_pointer == 90 && y_pointer == 37)
||(x_pointer == 91 && y_pointer == 37)
||(x_pointer == 92 && y_pointer == 37)
||(x_pointer == 93 && y_pointer == 37)
||(x_pointer == 94 && y_pointer == 37)
||(x_pointer == 95 && y_pointer == 37)
||(x_pointer == 96 && y_pointer == 37)
||(x_pointer == 97 && y_pointer == 37)
||(x_pointer == 98 && y_pointer == 37)
||(x_pointer == 99 && y_pointer == 37)
||(x_pointer == 100 && y_pointer == 37)
||(x_pointer == 101 && y_pointer == 37)
||(x_pointer == 102 && y_pointer == 37)
||(x_pointer == 103 && y_pointer == 37)
||(x_pointer == 104 && y_pointer == 37)
||(x_pointer == 105 && y_pointer == 37)
||(x_pointer == 106 && y_pointer == 37)
||(x_pointer == 107 && y_pointer == 37)
||(x_pointer == 108 && y_pointer == 37)
||(x_pointer == 109 && y_pointer == 37)
||(x_pointer == 110 && y_pointer == 37)
||(x_pointer == 111 && y_pointer == 37)
||(x_pointer == 112 && y_pointer == 37)
||(x_pointer == 155 && y_pointer == 37)
||(x_pointer == 156 && y_pointer == 37)
||(x_pointer == 157 && y_pointer == 37)
||(x_pointer == 2 && y_pointer == 38)
||(x_pointer == 3 && y_pointer == 38)
||(x_pointer == 4 && y_pointer == 38)
||(x_pointer == 50 && y_pointer == 38)
||(x_pointer == 51 && y_pointer == 38)
||(x_pointer == 52 && y_pointer == 38)
||(x_pointer == 53 && y_pointer == 38)
||(x_pointer == 54 && y_pointer == 38)
||(x_pointer == 55 && y_pointer == 38)
||(x_pointer == 56 && y_pointer == 38)
||(x_pointer == 57 && y_pointer == 38)
||(x_pointer == 58 && y_pointer == 38)
||(x_pointer == 59 && y_pointer == 38)
||(x_pointer == 60 && y_pointer == 38)
||(x_pointer == 61 && y_pointer == 38)
||(x_pointer == 62 && y_pointer == 38)
||(x_pointer == 63 && y_pointer == 38)
||(x_pointer == 64 && y_pointer == 38)
||(x_pointer == 65 && y_pointer == 38)
||(x_pointer == 66 && y_pointer == 38)
||(x_pointer == 67 && y_pointer == 38)
||(x_pointer == 68 && y_pointer == 38)
||(x_pointer == 69 && y_pointer == 38)
||(x_pointer == 70 && y_pointer == 38)
||(x_pointer == 71 && y_pointer == 38)
||(x_pointer == 72 && y_pointer == 38)
||(x_pointer == 73 && y_pointer == 38)
||(x_pointer == 89 && y_pointer == 38)
||(x_pointer == 90 && y_pointer == 38)
||(x_pointer == 91 && y_pointer == 38)
||(x_pointer == 92 && y_pointer == 38)
||(x_pointer == 93 && y_pointer == 38)
||(x_pointer == 94 && y_pointer == 38)
||(x_pointer == 95 && y_pointer == 38)
||(x_pointer == 96 && y_pointer == 38)
||(x_pointer == 97 && y_pointer == 38)
||(x_pointer == 98 && y_pointer == 38)
||(x_pointer == 99 && y_pointer == 38)
||(x_pointer == 100 && y_pointer == 38)
||(x_pointer == 101 && y_pointer == 38)
||(x_pointer == 102 && y_pointer == 38)
||(x_pointer == 103 && y_pointer == 38)
||(x_pointer == 104 && y_pointer == 38)
||(x_pointer == 105 && y_pointer == 38)
||(x_pointer == 106 && y_pointer == 38)
||(x_pointer == 107 && y_pointer == 38)
||(x_pointer == 108 && y_pointer == 38)
||(x_pointer == 109 && y_pointer == 38)
||(x_pointer == 110 && y_pointer == 38)
||(x_pointer == 111 && y_pointer == 38)
||(x_pointer == 112 && y_pointer == 38)
||(x_pointer == 155 && y_pointer == 38)
||(x_pointer == 156 && y_pointer == 38)
||(x_pointer == 157 && y_pointer == 38)
||(x_pointer == 2 && y_pointer == 39)
||(x_pointer == 3 && y_pointer == 39)
||(x_pointer == 4 && y_pointer == 39)
||(x_pointer == 50 && y_pointer == 39)
||(x_pointer == 51 && y_pointer == 39)
||(x_pointer == 52 && y_pointer == 39)
||(x_pointer == 53 && y_pointer == 39)
||(x_pointer == 54 && y_pointer == 39)
||(x_pointer == 55 && y_pointer == 39)
||(x_pointer == 56 && y_pointer == 39)
||(x_pointer == 57 && y_pointer == 39)
||(x_pointer == 58 && y_pointer == 39)
||(x_pointer == 59 && y_pointer == 39)
||(x_pointer == 60 && y_pointer == 39)
||(x_pointer == 61 && y_pointer == 39)
||(x_pointer == 62 && y_pointer == 39)
||(x_pointer == 63 && y_pointer == 39)
||(x_pointer == 64 && y_pointer == 39)
||(x_pointer == 65 && y_pointer == 39)
||(x_pointer == 66 && y_pointer == 39)
||(x_pointer == 67 && y_pointer == 39)
||(x_pointer == 68 && y_pointer == 39)
||(x_pointer == 69 && y_pointer == 39)
||(x_pointer == 70 && y_pointer == 39)
||(x_pointer == 71 && y_pointer == 39)
||(x_pointer == 72 && y_pointer == 39)
||(x_pointer == 73 && y_pointer == 39)
||(x_pointer == 89 && y_pointer == 39)
||(x_pointer == 90 && y_pointer == 39)
||(x_pointer == 91 && y_pointer == 39)
||(x_pointer == 92 && y_pointer == 39)
||(x_pointer == 93 && y_pointer == 39)
||(x_pointer == 94 && y_pointer == 39)
||(x_pointer == 95 && y_pointer == 39)
||(x_pointer == 96 && y_pointer == 39)
||(x_pointer == 97 && y_pointer == 39)
||(x_pointer == 98 && y_pointer == 39)
||(x_pointer == 99 && y_pointer == 39)
||(x_pointer == 100 && y_pointer == 39)
||(x_pointer == 101 && y_pointer == 39)
||(x_pointer == 102 && y_pointer == 39)
||(x_pointer == 103 && y_pointer == 39)
||(x_pointer == 104 && y_pointer == 39)
||(x_pointer == 105 && y_pointer == 39)
||(x_pointer == 106 && y_pointer == 39)
||(x_pointer == 107 && y_pointer == 39)
||(x_pointer == 108 && y_pointer == 39)
||(x_pointer == 109 && y_pointer == 39)
||(x_pointer == 110 && y_pointer == 39)
||(x_pointer == 111 && y_pointer == 39)
||(x_pointer == 112 && y_pointer == 39)
||(x_pointer == 155 && y_pointer == 39)
||(x_pointer == 156 && y_pointer == 39)
||(x_pointer == 157 && y_pointer == 39)
||(x_pointer == 2 && y_pointer == 40)
||(x_pointer == 3 && y_pointer == 40)
||(x_pointer == 4 && y_pointer == 40)
||(x_pointer == 50 && y_pointer == 40)
||(x_pointer == 51 && y_pointer == 40)
||(x_pointer == 52 && y_pointer == 40)
||(x_pointer == 53 && y_pointer == 40)
||(x_pointer == 54 && y_pointer == 40)
||(x_pointer == 55 && y_pointer == 40)
||(x_pointer == 56 && y_pointer == 40)
||(x_pointer == 57 && y_pointer == 40)
||(x_pointer == 58 && y_pointer == 40)
||(x_pointer == 59 && y_pointer == 40)
||(x_pointer == 60 && y_pointer == 40)
||(x_pointer == 61 && y_pointer == 40)
||(x_pointer == 62 && y_pointer == 40)
||(x_pointer == 63 && y_pointer == 40)
||(x_pointer == 64 && y_pointer == 40)
||(x_pointer == 65 && y_pointer == 40)
||(x_pointer == 66 && y_pointer == 40)
||(x_pointer == 67 && y_pointer == 40)
||(x_pointer == 68 && y_pointer == 40)
||(x_pointer == 69 && y_pointer == 40)
||(x_pointer == 70 && y_pointer == 40)
||(x_pointer == 71 && y_pointer == 40)
||(x_pointer == 72 && y_pointer == 40)
||(x_pointer == 73 && y_pointer == 40)
||(x_pointer == 89 && y_pointer == 40)
||(x_pointer == 90 && y_pointer == 40)
||(x_pointer == 91 && y_pointer == 40)
||(x_pointer == 92 && y_pointer == 40)
||(x_pointer == 93 && y_pointer == 40)
||(x_pointer == 94 && y_pointer == 40)
||(x_pointer == 95 && y_pointer == 40)
||(x_pointer == 96 && y_pointer == 40)
||(x_pointer == 97 && y_pointer == 40)
||(x_pointer == 98 && y_pointer == 40)
||(x_pointer == 99 && y_pointer == 40)
||(x_pointer == 100 && y_pointer == 40)
||(x_pointer == 101 && y_pointer == 40)
||(x_pointer == 102 && y_pointer == 40)
||(x_pointer == 103 && y_pointer == 40)
||(x_pointer == 104 && y_pointer == 40)
||(x_pointer == 105 && y_pointer == 40)
||(x_pointer == 106 && y_pointer == 40)
||(x_pointer == 107 && y_pointer == 40)
||(x_pointer == 108 && y_pointer == 40)
||(x_pointer == 109 && y_pointer == 40)
||(x_pointer == 110 && y_pointer == 40)
||(x_pointer == 111 && y_pointer == 40)
||(x_pointer == 112 && y_pointer == 40)
||(x_pointer == 155 && y_pointer == 40)
||(x_pointer == 156 && y_pointer == 40)
||(x_pointer == 157 && y_pointer == 40)
||(x_pointer == 2 && y_pointer == 41)
||(x_pointer == 3 && y_pointer == 41)
||(x_pointer == 4 && y_pointer == 41)
||(x_pointer == 50 && y_pointer == 41)
||(x_pointer == 51 && y_pointer == 41)
||(x_pointer == 52 && y_pointer == 41)
||(x_pointer == 53 && y_pointer == 41)
||(x_pointer == 54 && y_pointer == 41)
||(x_pointer == 55 && y_pointer == 41)
||(x_pointer == 56 && y_pointer == 41)
||(x_pointer == 57 && y_pointer == 41)
||(x_pointer == 58 && y_pointer == 41)
||(x_pointer == 59 && y_pointer == 41)
||(x_pointer == 60 && y_pointer == 41)
||(x_pointer == 61 && y_pointer == 41)
||(x_pointer == 62 && y_pointer == 41)
||(x_pointer == 63 && y_pointer == 41)
||(x_pointer == 64 && y_pointer == 41)
||(x_pointer == 65 && y_pointer == 41)
||(x_pointer == 66 && y_pointer == 41)
||(x_pointer == 67 && y_pointer == 41)
||(x_pointer == 68 && y_pointer == 41)
||(x_pointer == 69 && y_pointer == 41)
||(x_pointer == 70 && y_pointer == 41)
||(x_pointer == 71 && y_pointer == 41)
||(x_pointer == 72 && y_pointer == 41)
||(x_pointer == 73 && y_pointer == 41)
||(x_pointer == 89 && y_pointer == 41)
||(x_pointer == 90 && y_pointer == 41)
||(x_pointer == 91 && y_pointer == 41)
||(x_pointer == 92 && y_pointer == 41)
||(x_pointer == 93 && y_pointer == 41)
||(x_pointer == 94 && y_pointer == 41)
||(x_pointer == 95 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 99 && y_pointer == 41)
||(x_pointer == 100 && y_pointer == 41)
||(x_pointer == 101 && y_pointer == 41)
||(x_pointer == 102 && y_pointer == 41)
||(x_pointer == 103 && y_pointer == 41)
||(x_pointer == 104 && y_pointer == 41)
||(x_pointer == 105 && y_pointer == 41)
||(x_pointer == 106 && y_pointer == 41)
||(x_pointer == 107 && y_pointer == 41)
||(x_pointer == 108 && y_pointer == 41)
||(x_pointer == 109 && y_pointer == 41)
||(x_pointer == 110 && y_pointer == 41)
||(x_pointer == 111 && y_pointer == 41)
||(x_pointer == 112 && y_pointer == 41)
||(x_pointer == 155 && y_pointer == 41)
||(x_pointer == 156 && y_pointer == 41)
||(x_pointer == 157 && y_pointer == 41)
||(x_pointer == 2 && y_pointer == 42)
||(x_pointer == 3 && y_pointer == 42)
||(x_pointer == 4 && y_pointer == 42)
||(x_pointer == 50 && y_pointer == 42)
||(x_pointer == 51 && y_pointer == 42)
||(x_pointer == 52 && y_pointer == 42)
||(x_pointer == 53 && y_pointer == 42)
||(x_pointer == 54 && y_pointer == 42)
||(x_pointer == 55 && y_pointer == 42)
||(x_pointer == 56 && y_pointer == 42)
||(x_pointer == 57 && y_pointer == 42)
||(x_pointer == 58 && y_pointer == 42)
||(x_pointer == 59 && y_pointer == 42)
||(x_pointer == 60 && y_pointer == 42)
||(x_pointer == 61 && y_pointer == 42)
||(x_pointer == 62 && y_pointer == 42)
||(x_pointer == 63 && y_pointer == 42)
||(x_pointer == 64 && y_pointer == 42)
||(x_pointer == 65 && y_pointer == 42)
||(x_pointer == 66 && y_pointer == 42)
||(x_pointer == 67 && y_pointer == 42)
||(x_pointer == 68 && y_pointer == 42)
||(x_pointer == 69 && y_pointer == 42)
||(x_pointer == 70 && y_pointer == 42)
||(x_pointer == 71 && y_pointer == 42)
||(x_pointer == 72 && y_pointer == 42)
||(x_pointer == 73 && y_pointer == 42)
||(x_pointer == 89 && y_pointer == 42)
||(x_pointer == 90 && y_pointer == 42)
||(x_pointer == 91 && y_pointer == 42)
||(x_pointer == 92 && y_pointer == 42)
||(x_pointer == 93 && y_pointer == 42)
||(x_pointer == 94 && y_pointer == 42)
||(x_pointer == 95 && y_pointer == 42)
||(x_pointer == 96 && y_pointer == 42)
||(x_pointer == 97 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 99 && y_pointer == 42)
||(x_pointer == 100 && y_pointer == 42)
||(x_pointer == 101 && y_pointer == 42)
||(x_pointer == 102 && y_pointer == 42)
||(x_pointer == 103 && y_pointer == 42)
||(x_pointer == 104 && y_pointer == 42)
||(x_pointer == 105 && y_pointer == 42)
||(x_pointer == 106 && y_pointer == 42)
||(x_pointer == 107 && y_pointer == 42)
||(x_pointer == 108 && y_pointer == 42)
||(x_pointer == 109 && y_pointer == 42)
||(x_pointer == 110 && y_pointer == 42)
||(x_pointer == 111 && y_pointer == 42)
||(x_pointer == 112 && y_pointer == 42)
||(x_pointer == 155 && y_pointer == 42)
||(x_pointer == 156 && y_pointer == 42)
||(x_pointer == 157 && y_pointer == 42)
||(x_pointer == 2 && y_pointer == 43)
||(x_pointer == 3 && y_pointer == 43)
||(x_pointer == 4 && y_pointer == 43)
||(x_pointer == 50 && y_pointer == 43)
||(x_pointer == 51 && y_pointer == 43)
||(x_pointer == 52 && y_pointer == 43)
||(x_pointer == 53 && y_pointer == 43)
||(x_pointer == 54 && y_pointer == 43)
||(x_pointer == 55 && y_pointer == 43)
||(x_pointer == 56 && y_pointer == 43)
||(x_pointer == 57 && y_pointer == 43)
||(x_pointer == 58 && y_pointer == 43)
||(x_pointer == 59 && y_pointer == 43)
||(x_pointer == 60 && y_pointer == 43)
||(x_pointer == 61 && y_pointer == 43)
||(x_pointer == 62 && y_pointer == 43)
||(x_pointer == 63 && y_pointer == 43)
||(x_pointer == 64 && y_pointer == 43)
||(x_pointer == 65 && y_pointer == 43)
||(x_pointer == 66 && y_pointer == 43)
||(x_pointer == 67 && y_pointer == 43)
||(x_pointer == 68 && y_pointer == 43)
||(x_pointer == 69 && y_pointer == 43)
||(x_pointer == 70 && y_pointer == 43)
||(x_pointer == 71 && y_pointer == 43)
||(x_pointer == 72 && y_pointer == 43)
||(x_pointer == 73 && y_pointer == 43)
||(x_pointer == 89 && y_pointer == 43)
||(x_pointer == 90 && y_pointer == 43)
||(x_pointer == 91 && y_pointer == 43)
||(x_pointer == 92 && y_pointer == 43)
||(x_pointer == 93 && y_pointer == 43)
||(x_pointer == 94 && y_pointer == 43)
||(x_pointer == 95 && y_pointer == 43)
||(x_pointer == 96 && y_pointer == 43)
||(x_pointer == 97 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 99 && y_pointer == 43)
||(x_pointer == 100 && y_pointer == 43)
||(x_pointer == 101 && y_pointer == 43)
||(x_pointer == 102 && y_pointer == 43)
||(x_pointer == 103 && y_pointer == 43)
||(x_pointer == 104 && y_pointer == 43)
||(x_pointer == 105 && y_pointer == 43)
||(x_pointer == 106 && y_pointer == 43)
||(x_pointer == 107 && y_pointer == 43)
||(x_pointer == 108 && y_pointer == 43)
||(x_pointer == 109 && y_pointer == 43)
||(x_pointer == 110 && y_pointer == 43)
||(x_pointer == 111 && y_pointer == 43)
||(x_pointer == 112 && y_pointer == 43)
||(x_pointer == 155 && y_pointer == 43)
||(x_pointer == 156 && y_pointer == 43)
||(x_pointer == 157 && y_pointer == 43)
||(x_pointer == 2 && y_pointer == 44)
||(x_pointer == 3 && y_pointer == 44)
||(x_pointer == 4 && y_pointer == 44)
||(x_pointer == 50 && y_pointer == 44)
||(x_pointer == 51 && y_pointer == 44)
||(x_pointer == 52 && y_pointer == 44)
||(x_pointer == 53 && y_pointer == 44)
||(x_pointer == 54 && y_pointer == 44)
||(x_pointer == 55 && y_pointer == 44)
||(x_pointer == 56 && y_pointer == 44)
||(x_pointer == 57 && y_pointer == 44)
||(x_pointer == 58 && y_pointer == 44)
||(x_pointer == 59 && y_pointer == 44)
||(x_pointer == 60 && y_pointer == 44)
||(x_pointer == 61 && y_pointer == 44)
||(x_pointer == 62 && y_pointer == 44)
||(x_pointer == 63 && y_pointer == 44)
||(x_pointer == 64 && y_pointer == 44)
||(x_pointer == 65 && y_pointer == 44)
||(x_pointer == 66 && y_pointer == 44)
||(x_pointer == 67 && y_pointer == 44)
||(x_pointer == 68 && y_pointer == 44)
||(x_pointer == 69 && y_pointer == 44)
||(x_pointer == 70 && y_pointer == 44)
||(x_pointer == 71 && y_pointer == 44)
||(x_pointer == 72 && y_pointer == 44)
||(x_pointer == 73 && y_pointer == 44)
||(x_pointer == 89 && y_pointer == 44)
||(x_pointer == 90 && y_pointer == 44)
||(x_pointer == 91 && y_pointer == 44)
||(x_pointer == 92 && y_pointer == 44)
||(x_pointer == 93 && y_pointer == 44)
||(x_pointer == 94 && y_pointer == 44)
||(x_pointer == 95 && y_pointer == 44)
||(x_pointer == 96 && y_pointer == 44)
||(x_pointer == 97 && y_pointer == 44)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 99 && y_pointer == 44)
||(x_pointer == 100 && y_pointer == 44)
||(x_pointer == 101 && y_pointer == 44)
||(x_pointer == 102 && y_pointer == 44)
||(x_pointer == 103 && y_pointer == 44)
||(x_pointer == 104 && y_pointer == 44)
||(x_pointer == 105 && y_pointer == 44)
||(x_pointer == 106 && y_pointer == 44)
||(x_pointer == 107 && y_pointer == 44)
||(x_pointer == 108 && y_pointer == 44)
||(x_pointer == 109 && y_pointer == 44)
||(x_pointer == 110 && y_pointer == 44)
||(x_pointer == 111 && y_pointer == 44)
||(x_pointer == 112 && y_pointer == 44)
||(x_pointer == 155 && y_pointer == 44)
||(x_pointer == 156 && y_pointer == 44)
||(x_pointer == 157 && y_pointer == 44)
||(x_pointer == 2 && y_pointer == 45)
||(x_pointer == 3 && y_pointer == 45)
||(x_pointer == 4 && y_pointer == 45)
||(x_pointer == 50 && y_pointer == 45)
||(x_pointer == 51 && y_pointer == 45)
||(x_pointer == 52 && y_pointer == 45)
||(x_pointer == 53 && y_pointer == 45)
||(x_pointer == 54 && y_pointer == 45)
||(x_pointer == 55 && y_pointer == 45)
||(x_pointer == 56 && y_pointer == 45)
||(x_pointer == 57 && y_pointer == 45)
||(x_pointer == 58 && y_pointer == 45)
||(x_pointer == 59 && y_pointer == 45)
||(x_pointer == 60 && y_pointer == 45)
||(x_pointer == 61 && y_pointer == 45)
||(x_pointer == 62 && y_pointer == 45)
||(x_pointer == 63 && y_pointer == 45)
||(x_pointer == 64 && y_pointer == 45)
||(x_pointer == 65 && y_pointer == 45)
||(x_pointer == 66 && y_pointer == 45)
||(x_pointer == 67 && y_pointer == 45)
||(x_pointer == 68 && y_pointer == 45)
||(x_pointer == 69 && y_pointer == 45)
||(x_pointer == 70 && y_pointer == 45)
||(x_pointer == 71 && y_pointer == 45)
||(x_pointer == 72 && y_pointer == 45)
||(x_pointer == 73 && y_pointer == 45)
||(x_pointer == 89 && y_pointer == 45)
||(x_pointer == 90 && y_pointer == 45)
||(x_pointer == 91 && y_pointer == 45)
||(x_pointer == 92 && y_pointer == 45)
||(x_pointer == 93 && y_pointer == 45)
||(x_pointer == 94 && y_pointer == 45)
||(x_pointer == 95 && y_pointer == 45)
||(x_pointer == 96 && y_pointer == 45)
||(x_pointer == 97 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 99 && y_pointer == 45)
||(x_pointer == 100 && y_pointer == 45)
||(x_pointer == 101 && y_pointer == 45)
||(x_pointer == 102 && y_pointer == 45)
||(x_pointer == 103 && y_pointer == 45)
||(x_pointer == 104 && y_pointer == 45)
||(x_pointer == 105 && y_pointer == 45)
||(x_pointer == 106 && y_pointer == 45)
||(x_pointer == 107 && y_pointer == 45)
||(x_pointer == 108 && y_pointer == 45)
||(x_pointer == 109 && y_pointer == 45)
||(x_pointer == 110 && y_pointer == 45)
||(x_pointer == 111 && y_pointer == 45)
||(x_pointer == 112 && y_pointer == 45)
||(x_pointer == 155 && y_pointer == 45)
||(x_pointer == 156 && y_pointer == 45)
||(x_pointer == 157 && y_pointer == 45)
||(x_pointer == 2 && y_pointer == 46)
||(x_pointer == 3 && y_pointer == 46)
||(x_pointer == 4 && y_pointer == 46)
||(x_pointer == 50 && y_pointer == 46)
||(x_pointer == 51 && y_pointer == 46)
||(x_pointer == 52 && y_pointer == 46)
||(x_pointer == 53 && y_pointer == 46)
||(x_pointer == 54 && y_pointer == 46)
||(x_pointer == 55 && y_pointer == 46)
||(x_pointer == 56 && y_pointer == 46)
||(x_pointer == 57 && y_pointer == 46)
||(x_pointer == 58 && y_pointer == 46)
||(x_pointer == 59 && y_pointer == 46)
||(x_pointer == 60 && y_pointer == 46)
||(x_pointer == 61 && y_pointer == 46)
||(x_pointer == 62 && y_pointer == 46)
||(x_pointer == 63 && y_pointer == 46)
||(x_pointer == 64 && y_pointer == 46)
||(x_pointer == 65 && y_pointer == 46)
||(x_pointer == 66 && y_pointer == 46)
||(x_pointer == 67 && y_pointer == 46)
||(x_pointer == 68 && y_pointer == 46)
||(x_pointer == 69 && y_pointer == 46)
||(x_pointer == 70 && y_pointer == 46)
||(x_pointer == 71 && y_pointer == 46)
||(x_pointer == 72 && y_pointer == 46)
||(x_pointer == 73 && y_pointer == 46)
||(x_pointer == 89 && y_pointer == 46)
||(x_pointer == 90 && y_pointer == 46)
||(x_pointer == 91 && y_pointer == 46)
||(x_pointer == 92 && y_pointer == 46)
||(x_pointer == 93 && y_pointer == 46)
||(x_pointer == 94 && y_pointer == 46)
||(x_pointer == 95 && y_pointer == 46)
||(x_pointer == 96 && y_pointer == 46)
||(x_pointer == 97 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 99 && y_pointer == 46)
||(x_pointer == 100 && y_pointer == 46)
||(x_pointer == 101 && y_pointer == 46)
||(x_pointer == 102 && y_pointer == 46)
||(x_pointer == 103 && y_pointer == 46)
||(x_pointer == 104 && y_pointer == 46)
||(x_pointer == 105 && y_pointer == 46)
||(x_pointer == 106 && y_pointer == 46)
||(x_pointer == 107 && y_pointer == 46)
||(x_pointer == 108 && y_pointer == 46)
||(x_pointer == 109 && y_pointer == 46)
||(x_pointer == 110 && y_pointer == 46)
||(x_pointer == 111 && y_pointer == 46)
||(x_pointer == 112 && y_pointer == 46)
||(x_pointer == 155 && y_pointer == 46)
||(x_pointer == 156 && y_pointer == 46)
||(x_pointer == 157 && y_pointer == 46)
||(x_pointer == 2 && y_pointer == 47)
||(x_pointer == 3 && y_pointer == 47)
||(x_pointer == 4 && y_pointer == 47)
||(x_pointer == 50 && y_pointer == 47)
||(x_pointer == 51 && y_pointer == 47)
||(x_pointer == 52 && y_pointer == 47)
||(x_pointer == 53 && y_pointer == 47)
||(x_pointer == 54 && y_pointer == 47)
||(x_pointer == 55 && y_pointer == 47)
||(x_pointer == 56 && y_pointer == 47)
||(x_pointer == 57 && y_pointer == 47)
||(x_pointer == 58 && y_pointer == 47)
||(x_pointer == 59 && y_pointer == 47)
||(x_pointer == 60 && y_pointer == 47)
||(x_pointer == 61 && y_pointer == 47)
||(x_pointer == 62 && y_pointer == 47)
||(x_pointer == 63 && y_pointer == 47)
||(x_pointer == 64 && y_pointer == 47)
||(x_pointer == 65 && y_pointer == 47)
||(x_pointer == 66 && y_pointer == 47)
||(x_pointer == 67 && y_pointer == 47)
||(x_pointer == 68 && y_pointer == 47)
||(x_pointer == 69 && y_pointer == 47)
||(x_pointer == 70 && y_pointer == 47)
||(x_pointer == 71 && y_pointer == 47)
||(x_pointer == 72 && y_pointer == 47)
||(x_pointer == 73 && y_pointer == 47)
||(x_pointer == 74 && y_pointer == 47)
||(x_pointer == 75 && y_pointer == 47)
||(x_pointer == 76 && y_pointer == 47)
||(x_pointer == 77 && y_pointer == 47)
||(x_pointer == 78 && y_pointer == 47)
||(x_pointer == 79 && y_pointer == 47)
||(x_pointer == 80 && y_pointer == 47)
||(x_pointer == 81 && y_pointer == 47)
||(x_pointer == 82 && y_pointer == 47)
||(x_pointer == 83 && y_pointer == 47)
||(x_pointer == 84 && y_pointer == 47)
||(x_pointer == 85 && y_pointer == 47)
||(x_pointer == 86 && y_pointer == 47)
||(x_pointer == 87 && y_pointer == 47)
||(x_pointer == 88 && y_pointer == 47)
||(x_pointer == 89 && y_pointer == 47)
||(x_pointer == 90 && y_pointer == 47)
||(x_pointer == 91 && y_pointer == 47)
||(x_pointer == 92 && y_pointer == 47)
||(x_pointer == 93 && y_pointer == 47)
||(x_pointer == 94 && y_pointer == 47)
||(x_pointer == 95 && y_pointer == 47)
||(x_pointer == 96 && y_pointer == 47)
||(x_pointer == 97 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 99 && y_pointer == 47)
||(x_pointer == 100 && y_pointer == 47)
||(x_pointer == 101 && y_pointer == 47)
||(x_pointer == 102 && y_pointer == 47)
||(x_pointer == 103 && y_pointer == 47)
||(x_pointer == 104 && y_pointer == 47)
||(x_pointer == 105 && y_pointer == 47)
||(x_pointer == 106 && y_pointer == 47)
||(x_pointer == 107 && y_pointer == 47)
||(x_pointer == 108 && y_pointer == 47)
||(x_pointer == 109 && y_pointer == 47)
||(x_pointer == 110 && y_pointer == 47)
||(x_pointer == 111 && y_pointer == 47)
||(x_pointer == 112 && y_pointer == 47)
||(x_pointer == 155 && y_pointer == 47)
||(x_pointer == 156 && y_pointer == 47)
||(x_pointer == 157 && y_pointer == 47)
||(x_pointer == 2 && y_pointer == 48)
||(x_pointer == 3 && y_pointer == 48)
||(x_pointer == 4 && y_pointer == 48)
||(x_pointer == 50 && y_pointer == 48)
||(x_pointer == 51 && y_pointer == 48)
||(x_pointer == 52 && y_pointer == 48)
||(x_pointer == 53 && y_pointer == 48)
||(x_pointer == 54 && y_pointer == 48)
||(x_pointer == 55 && y_pointer == 48)
||(x_pointer == 56 && y_pointer == 48)
||(x_pointer == 57 && y_pointer == 48)
||(x_pointer == 58 && y_pointer == 48)
||(x_pointer == 59 && y_pointer == 48)
||(x_pointer == 60 && y_pointer == 48)
||(x_pointer == 61 && y_pointer == 48)
||(x_pointer == 62 && y_pointer == 48)
||(x_pointer == 63 && y_pointer == 48)
||(x_pointer == 64 && y_pointer == 48)
||(x_pointer == 65 && y_pointer == 48)
||(x_pointer == 66 && y_pointer == 48)
||(x_pointer == 67 && y_pointer == 48)
||(x_pointer == 68 && y_pointer == 48)
||(x_pointer == 69 && y_pointer == 48)
||(x_pointer == 70 && y_pointer == 48)
||(x_pointer == 71 && y_pointer == 48)
||(x_pointer == 72 && y_pointer == 48)
||(x_pointer == 73 && y_pointer == 48)
||(x_pointer == 74 && y_pointer == 48)
||(x_pointer == 75 && y_pointer == 48)
||(x_pointer == 76 && y_pointer == 48)
||(x_pointer == 77 && y_pointer == 48)
||(x_pointer == 78 && y_pointer == 48)
||(x_pointer == 79 && y_pointer == 48)
||(x_pointer == 80 && y_pointer == 48)
||(x_pointer == 81 && y_pointer == 48)
||(x_pointer == 82 && y_pointer == 48)
||(x_pointer == 83 && y_pointer == 48)
||(x_pointer == 84 && y_pointer == 48)
||(x_pointer == 85 && y_pointer == 48)
||(x_pointer == 86 && y_pointer == 48)
||(x_pointer == 87 && y_pointer == 48)
||(x_pointer == 88 && y_pointer == 48)
||(x_pointer == 89 && y_pointer == 48)
||(x_pointer == 90 && y_pointer == 48)
||(x_pointer == 91 && y_pointer == 48)
||(x_pointer == 92 && y_pointer == 48)
||(x_pointer == 93 && y_pointer == 48)
||(x_pointer == 94 && y_pointer == 48)
||(x_pointer == 95 && y_pointer == 48)
||(x_pointer == 96 && y_pointer == 48)
||(x_pointer == 97 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 48)
||(x_pointer == 99 && y_pointer == 48)
||(x_pointer == 100 && y_pointer == 48)
||(x_pointer == 101 && y_pointer == 48)
||(x_pointer == 102 && y_pointer == 48)
||(x_pointer == 103 && y_pointer == 48)
||(x_pointer == 104 && y_pointer == 48)
||(x_pointer == 105 && y_pointer == 48)
||(x_pointer == 106 && y_pointer == 48)
||(x_pointer == 107 && y_pointer == 48)
||(x_pointer == 108 && y_pointer == 48)
||(x_pointer == 109 && y_pointer == 48)
||(x_pointer == 110 && y_pointer == 48)
||(x_pointer == 111 && y_pointer == 48)
||(x_pointer == 112 && y_pointer == 48)
||(x_pointer == 155 && y_pointer == 48)
||(x_pointer == 156 && y_pointer == 48)
||(x_pointer == 157 && y_pointer == 48)
||(x_pointer == 2 && y_pointer == 49)
||(x_pointer == 3 && y_pointer == 49)
||(x_pointer == 4 && y_pointer == 49)
||(x_pointer == 50 && y_pointer == 49)
||(x_pointer == 51 && y_pointer == 49)
||(x_pointer == 52 && y_pointer == 49)
||(x_pointer == 53 && y_pointer == 49)
||(x_pointer == 54 && y_pointer == 49)
||(x_pointer == 55 && y_pointer == 49)
||(x_pointer == 56 && y_pointer == 49)
||(x_pointer == 57 && y_pointer == 49)
||(x_pointer == 58 && y_pointer == 49)
||(x_pointer == 59 && y_pointer == 49)
||(x_pointer == 60 && y_pointer == 49)
||(x_pointer == 61 && y_pointer == 49)
||(x_pointer == 62 && y_pointer == 49)
||(x_pointer == 63 && y_pointer == 49)
||(x_pointer == 64 && y_pointer == 49)
||(x_pointer == 65 && y_pointer == 49)
||(x_pointer == 66 && y_pointer == 49)
||(x_pointer == 67 && y_pointer == 49)
||(x_pointer == 68 && y_pointer == 49)
||(x_pointer == 69 && y_pointer == 49)
||(x_pointer == 70 && y_pointer == 49)
||(x_pointer == 71 && y_pointer == 49)
||(x_pointer == 72 && y_pointer == 49)
||(x_pointer == 73 && y_pointer == 49)
||(x_pointer == 74 && y_pointer == 49)
||(x_pointer == 75 && y_pointer == 49)
||(x_pointer == 76 && y_pointer == 49)
||(x_pointer == 77 && y_pointer == 49)
||(x_pointer == 78 && y_pointer == 49)
||(x_pointer == 79 && y_pointer == 49)
||(x_pointer == 80 && y_pointer == 49)
||(x_pointer == 81 && y_pointer == 49)
||(x_pointer == 82 && y_pointer == 49)
||(x_pointer == 83 && y_pointer == 49)
||(x_pointer == 84 && y_pointer == 49)
||(x_pointer == 85 && y_pointer == 49)
||(x_pointer == 86 && y_pointer == 49)
||(x_pointer == 87 && y_pointer == 49)
||(x_pointer == 88 && y_pointer == 49)
||(x_pointer == 89 && y_pointer == 49)
||(x_pointer == 90 && y_pointer == 49)
||(x_pointer == 91 && y_pointer == 49)
||(x_pointer == 92 && y_pointer == 49)
||(x_pointer == 93 && y_pointer == 49)
||(x_pointer == 94 && y_pointer == 49)
||(x_pointer == 95 && y_pointer == 49)
||(x_pointer == 96 && y_pointer == 49)
||(x_pointer == 97 && y_pointer == 49)
||(x_pointer == 98 && y_pointer == 49)
||(x_pointer == 99 && y_pointer == 49)
||(x_pointer == 100 && y_pointer == 49)
||(x_pointer == 101 && y_pointer == 49)
||(x_pointer == 102 && y_pointer == 49)
||(x_pointer == 103 && y_pointer == 49)
||(x_pointer == 104 && y_pointer == 49)
||(x_pointer == 105 && y_pointer == 49)
||(x_pointer == 106 && y_pointer == 49)
||(x_pointer == 107 && y_pointer == 49)
||(x_pointer == 108 && y_pointer == 49)
||(x_pointer == 109 && y_pointer == 49)
||(x_pointer == 110 && y_pointer == 49)
||(x_pointer == 111 && y_pointer == 49)
||(x_pointer == 112 && y_pointer == 49)
||(x_pointer == 155 && y_pointer == 49)
||(x_pointer == 156 && y_pointer == 49)
||(x_pointer == 157 && y_pointer == 49)
||(x_pointer == 2 && y_pointer == 50)
||(x_pointer == 3 && y_pointer == 50)
||(x_pointer == 4 && y_pointer == 50)
||(x_pointer == 71 && y_pointer == 50)
||(x_pointer == 72 && y_pointer == 50)
||(x_pointer == 73 && y_pointer == 50)
||(x_pointer == 74 && y_pointer == 50)
||(x_pointer == 75 && y_pointer == 50)
||(x_pointer == 76 && y_pointer == 50)
||(x_pointer == 77 && y_pointer == 50)
||(x_pointer == 78 && y_pointer == 50)
||(x_pointer == 79 && y_pointer == 50)
||(x_pointer == 80 && y_pointer == 50)
||(x_pointer == 81 && y_pointer == 50)
||(x_pointer == 82 && y_pointer == 50)
||(x_pointer == 83 && y_pointer == 50)
||(x_pointer == 84 && y_pointer == 50)
||(x_pointer == 85 && y_pointer == 50)
||(x_pointer == 86 && y_pointer == 50)
||(x_pointer == 87 && y_pointer == 50)
||(x_pointer == 88 && y_pointer == 50)
||(x_pointer == 89 && y_pointer == 50)
||(x_pointer == 90 && y_pointer == 50)
||(x_pointer == 91 && y_pointer == 50)
||(x_pointer == 155 && y_pointer == 50)
||(x_pointer == 156 && y_pointer == 50)
||(x_pointer == 157 && y_pointer == 50)
||(x_pointer == 2 && y_pointer == 51)
||(x_pointer == 3 && y_pointer == 51)
||(x_pointer == 4 && y_pointer == 51)
||(x_pointer == 71 && y_pointer == 51)
||(x_pointer == 72 && y_pointer == 51)
||(x_pointer == 73 && y_pointer == 51)
||(x_pointer == 74 && y_pointer == 51)
||(x_pointer == 75 && y_pointer == 51)
||(x_pointer == 76 && y_pointer == 51)
||(x_pointer == 77 && y_pointer == 51)
||(x_pointer == 78 && y_pointer == 51)
||(x_pointer == 79 && y_pointer == 51)
||(x_pointer == 80 && y_pointer == 51)
||(x_pointer == 81 && y_pointer == 51)
||(x_pointer == 82 && y_pointer == 51)
||(x_pointer == 83 && y_pointer == 51)
||(x_pointer == 84 && y_pointer == 51)
||(x_pointer == 85 && y_pointer == 51)
||(x_pointer == 86 && y_pointer == 51)
||(x_pointer == 87 && y_pointer == 51)
||(x_pointer == 88 && y_pointer == 51)
||(x_pointer == 89 && y_pointer == 51)
||(x_pointer == 90 && y_pointer == 51)
||(x_pointer == 91 && y_pointer == 51)
||(x_pointer == 155 && y_pointer == 51)
||(x_pointer == 156 && y_pointer == 51)
||(x_pointer == 157 && y_pointer == 51)
||(x_pointer == 2 && y_pointer == 52)
||(x_pointer == 3 && y_pointer == 52)
||(x_pointer == 4 && y_pointer == 52)
||(x_pointer == 71 && y_pointer == 52)
||(x_pointer == 72 && y_pointer == 52)
||(x_pointer == 73 && y_pointer == 52)
||(x_pointer == 74 && y_pointer == 52)
||(x_pointer == 75 && y_pointer == 52)
||(x_pointer == 76 && y_pointer == 52)
||(x_pointer == 77 && y_pointer == 52)
||(x_pointer == 78 && y_pointer == 52)
||(x_pointer == 79 && y_pointer == 52)
||(x_pointer == 80 && y_pointer == 52)
||(x_pointer == 81 && y_pointer == 52)
||(x_pointer == 82 && y_pointer == 52)
||(x_pointer == 83 && y_pointer == 52)
||(x_pointer == 84 && y_pointer == 52)
||(x_pointer == 85 && y_pointer == 52)
||(x_pointer == 86 && y_pointer == 52)
||(x_pointer == 87 && y_pointer == 52)
||(x_pointer == 88 && y_pointer == 52)
||(x_pointer == 89 && y_pointer == 52)
||(x_pointer == 90 && y_pointer == 52)
||(x_pointer == 91 && y_pointer == 52)
||(x_pointer == 155 && y_pointer == 52)
||(x_pointer == 156 && y_pointer == 52)
||(x_pointer == 157 && y_pointer == 52)
||(x_pointer == 2 && y_pointer == 53)
||(x_pointer == 3 && y_pointer == 53)
||(x_pointer == 4 && y_pointer == 53)
||(x_pointer == 71 && y_pointer == 53)
||(x_pointer == 72 && y_pointer == 53)
||(x_pointer == 73 && y_pointer == 53)
||(x_pointer == 74 && y_pointer == 53)
||(x_pointer == 75 && y_pointer == 53)
||(x_pointer == 76 && y_pointer == 53)
||(x_pointer == 77 && y_pointer == 53)
||(x_pointer == 78 && y_pointer == 53)
||(x_pointer == 79 && y_pointer == 53)
||(x_pointer == 80 && y_pointer == 53)
||(x_pointer == 81 && y_pointer == 53)
||(x_pointer == 82 && y_pointer == 53)
||(x_pointer == 83 && y_pointer == 53)
||(x_pointer == 84 && y_pointer == 53)
||(x_pointer == 85 && y_pointer == 53)
||(x_pointer == 86 && y_pointer == 53)
||(x_pointer == 87 && y_pointer == 53)
||(x_pointer == 88 && y_pointer == 53)
||(x_pointer == 89 && y_pointer == 53)
||(x_pointer == 90 && y_pointer == 53)
||(x_pointer == 91 && y_pointer == 53)
||(x_pointer == 155 && y_pointer == 53)
||(x_pointer == 156 && y_pointer == 53)
||(x_pointer == 157 && y_pointer == 53)
||(x_pointer == 2 && y_pointer == 54)
||(x_pointer == 3 && y_pointer == 54)
||(x_pointer == 4 && y_pointer == 54)
||(x_pointer == 71 && y_pointer == 54)
||(x_pointer == 72 && y_pointer == 54)
||(x_pointer == 73 && y_pointer == 54)
||(x_pointer == 74 && y_pointer == 54)
||(x_pointer == 75 && y_pointer == 54)
||(x_pointer == 76 && y_pointer == 54)
||(x_pointer == 77 && y_pointer == 54)
||(x_pointer == 78 && y_pointer == 54)
||(x_pointer == 79 && y_pointer == 54)
||(x_pointer == 80 && y_pointer == 54)
||(x_pointer == 81 && y_pointer == 54)
||(x_pointer == 82 && y_pointer == 54)
||(x_pointer == 83 && y_pointer == 54)
||(x_pointer == 84 && y_pointer == 54)
||(x_pointer == 85 && y_pointer == 54)
||(x_pointer == 86 && y_pointer == 54)
||(x_pointer == 87 && y_pointer == 54)
||(x_pointer == 88 && y_pointer == 54)
||(x_pointer == 89 && y_pointer == 54)
||(x_pointer == 90 && y_pointer == 54)
||(x_pointer == 91 && y_pointer == 54)
||(x_pointer == 155 && y_pointer == 54)
||(x_pointer == 156 && y_pointer == 54)
||(x_pointer == 157 && y_pointer == 54)
||(x_pointer == 2 && y_pointer == 55)
||(x_pointer == 3 && y_pointer == 55)
||(x_pointer == 4 && y_pointer == 55)
||(x_pointer == 71 && y_pointer == 55)
||(x_pointer == 72 && y_pointer == 55)
||(x_pointer == 73 && y_pointer == 55)
||(x_pointer == 74 && y_pointer == 55)
||(x_pointer == 75 && y_pointer == 55)
||(x_pointer == 76 && y_pointer == 55)
||(x_pointer == 77 && y_pointer == 55)
||(x_pointer == 78 && y_pointer == 55)
||(x_pointer == 79 && y_pointer == 55)
||(x_pointer == 80 && y_pointer == 55)
||(x_pointer == 81 && y_pointer == 55)
||(x_pointer == 82 && y_pointer == 55)
||(x_pointer == 83 && y_pointer == 55)
||(x_pointer == 84 && y_pointer == 55)
||(x_pointer == 85 && y_pointer == 55)
||(x_pointer == 86 && y_pointer == 55)
||(x_pointer == 87 && y_pointer == 55)
||(x_pointer == 88 && y_pointer == 55)
||(x_pointer == 89 && y_pointer == 55)
||(x_pointer == 90 && y_pointer == 55)
||(x_pointer == 91 && y_pointer == 55)
||(x_pointer == 155 && y_pointer == 55)
||(x_pointer == 156 && y_pointer == 55)
||(x_pointer == 157 && y_pointer == 55)
||(x_pointer == 2 && y_pointer == 56)
||(x_pointer == 3 && y_pointer == 56)
||(x_pointer == 4 && y_pointer == 56)
||(x_pointer == 71 && y_pointer == 56)
||(x_pointer == 72 && y_pointer == 56)
||(x_pointer == 73 && y_pointer == 56)
||(x_pointer == 74 && y_pointer == 56)
||(x_pointer == 75 && y_pointer == 56)
||(x_pointer == 76 && y_pointer == 56)
||(x_pointer == 77 && y_pointer == 56)
||(x_pointer == 78 && y_pointer == 56)
||(x_pointer == 79 && y_pointer == 56)
||(x_pointer == 80 && y_pointer == 56)
||(x_pointer == 81 && y_pointer == 56)
||(x_pointer == 82 && y_pointer == 56)
||(x_pointer == 83 && y_pointer == 56)
||(x_pointer == 84 && y_pointer == 56)
||(x_pointer == 85 && y_pointer == 56)
||(x_pointer == 86 && y_pointer == 56)
||(x_pointer == 87 && y_pointer == 56)
||(x_pointer == 88 && y_pointer == 56)
||(x_pointer == 89 && y_pointer == 56)
||(x_pointer == 90 && y_pointer == 56)
||(x_pointer == 91 && y_pointer == 56)
||(x_pointer == 155 && y_pointer == 56)
||(x_pointer == 156 && y_pointer == 56)
||(x_pointer == 157 && y_pointer == 56)
||(x_pointer == 2 && y_pointer == 57)
||(x_pointer == 3 && y_pointer == 57)
||(x_pointer == 4 && y_pointer == 57)
||(x_pointer == 71 && y_pointer == 57)
||(x_pointer == 72 && y_pointer == 57)
||(x_pointer == 73 && y_pointer == 57)
||(x_pointer == 74 && y_pointer == 57)
||(x_pointer == 75 && y_pointer == 57)
||(x_pointer == 76 && y_pointer == 57)
||(x_pointer == 77 && y_pointer == 57)
||(x_pointer == 78 && y_pointer == 57)
||(x_pointer == 79 && y_pointer == 57)
||(x_pointer == 80 && y_pointer == 57)
||(x_pointer == 81 && y_pointer == 57)
||(x_pointer == 82 && y_pointer == 57)
||(x_pointer == 83 && y_pointer == 57)
||(x_pointer == 84 && y_pointer == 57)
||(x_pointer == 85 && y_pointer == 57)
||(x_pointer == 86 && y_pointer == 57)
||(x_pointer == 87 && y_pointer == 57)
||(x_pointer == 88 && y_pointer == 57)
||(x_pointer == 89 && y_pointer == 57)
||(x_pointer == 90 && y_pointer == 57)
||(x_pointer == 91 && y_pointer == 57)
||(x_pointer == 155 && y_pointer == 57)
||(x_pointer == 156 && y_pointer == 57)
||(x_pointer == 157 && y_pointer == 57)
||(x_pointer == 2 && y_pointer == 58)
||(x_pointer == 3 && y_pointer == 58)
||(x_pointer == 4 && y_pointer == 58)
||(x_pointer == 71 && y_pointer == 58)
||(x_pointer == 72 && y_pointer == 58)
||(x_pointer == 73 && y_pointer == 58)
||(x_pointer == 74 && y_pointer == 58)
||(x_pointer == 75 && y_pointer == 58)
||(x_pointer == 76 && y_pointer == 58)
||(x_pointer == 77 && y_pointer == 58)
||(x_pointer == 78 && y_pointer == 58)
||(x_pointer == 79 && y_pointer == 58)
||(x_pointer == 80 && y_pointer == 58)
||(x_pointer == 81 && y_pointer == 58)
||(x_pointer == 82 && y_pointer == 58)
||(x_pointer == 83 && y_pointer == 58)
||(x_pointer == 84 && y_pointer == 58)
||(x_pointer == 85 && y_pointer == 58)
||(x_pointer == 86 && y_pointer == 58)
||(x_pointer == 87 && y_pointer == 58)
||(x_pointer == 88 && y_pointer == 58)
||(x_pointer == 89 && y_pointer == 58)
||(x_pointer == 90 && y_pointer == 58)
||(x_pointer == 91 && y_pointer == 58)
||(x_pointer == 155 && y_pointer == 58)
||(x_pointer == 156 && y_pointer == 58)
||(x_pointer == 157 && y_pointer == 58)
||(x_pointer == 2 && y_pointer == 59)
||(x_pointer == 3 && y_pointer == 59)
||(x_pointer == 4 && y_pointer == 59)
||(x_pointer == 71 && y_pointer == 59)
||(x_pointer == 72 && y_pointer == 59)
||(x_pointer == 73 && y_pointer == 59)
||(x_pointer == 74 && y_pointer == 59)
||(x_pointer == 75 && y_pointer == 59)
||(x_pointer == 76 && y_pointer == 59)
||(x_pointer == 77 && y_pointer == 59)
||(x_pointer == 78 && y_pointer == 59)
||(x_pointer == 79 && y_pointer == 59)
||(x_pointer == 80 && y_pointer == 59)
||(x_pointer == 81 && y_pointer == 59)
||(x_pointer == 82 && y_pointer == 59)
||(x_pointer == 83 && y_pointer == 59)
||(x_pointer == 84 && y_pointer == 59)
||(x_pointer == 85 && y_pointer == 59)
||(x_pointer == 86 && y_pointer == 59)
||(x_pointer == 87 && y_pointer == 59)
||(x_pointer == 88 && y_pointer == 59)
||(x_pointer == 89 && y_pointer == 59)
||(x_pointer == 90 && y_pointer == 59)
||(x_pointer == 91 && y_pointer == 59)
||(x_pointer == 155 && y_pointer == 59)
||(x_pointer == 156 && y_pointer == 59)
||(x_pointer == 157 && y_pointer == 59)
||(x_pointer == 2 && y_pointer == 60)
||(x_pointer == 3 && y_pointer == 60)
||(x_pointer == 4 && y_pointer == 60)
||(x_pointer == 71 && y_pointer == 60)
||(x_pointer == 72 && y_pointer == 60)
||(x_pointer == 73 && y_pointer == 60)
||(x_pointer == 74 && y_pointer == 60)
||(x_pointer == 75 && y_pointer == 60)
||(x_pointer == 76 && y_pointer == 60)
||(x_pointer == 77 && y_pointer == 60)
||(x_pointer == 78 && y_pointer == 60)
||(x_pointer == 79 && y_pointer == 60)
||(x_pointer == 80 && y_pointer == 60)
||(x_pointer == 81 && y_pointer == 60)
||(x_pointer == 82 && y_pointer == 60)
||(x_pointer == 83 && y_pointer == 60)
||(x_pointer == 84 && y_pointer == 60)
||(x_pointer == 85 && y_pointer == 60)
||(x_pointer == 86 && y_pointer == 60)
||(x_pointer == 87 && y_pointer == 60)
||(x_pointer == 88 && y_pointer == 60)
||(x_pointer == 89 && y_pointer == 60)
||(x_pointer == 90 && y_pointer == 60)
||(x_pointer == 91 && y_pointer == 60)
||(x_pointer == 155 && y_pointer == 60)
||(x_pointer == 156 && y_pointer == 60)
||(x_pointer == 157 && y_pointer == 60)
||(x_pointer == 2 && y_pointer == 61)
||(x_pointer == 3 && y_pointer == 61)
||(x_pointer == 4 && y_pointer == 61)
||(x_pointer == 71 && y_pointer == 61)
||(x_pointer == 72 && y_pointer == 61)
||(x_pointer == 73 && y_pointer == 61)
||(x_pointer == 74 && y_pointer == 61)
||(x_pointer == 75 && y_pointer == 61)
||(x_pointer == 76 && y_pointer == 61)
||(x_pointer == 77 && y_pointer == 61)
||(x_pointer == 78 && y_pointer == 61)
||(x_pointer == 79 && y_pointer == 61)
||(x_pointer == 80 && y_pointer == 61)
||(x_pointer == 81 && y_pointer == 61)
||(x_pointer == 82 && y_pointer == 61)
||(x_pointer == 83 && y_pointer == 61)
||(x_pointer == 84 && y_pointer == 61)
||(x_pointer == 85 && y_pointer == 61)
||(x_pointer == 86 && y_pointer == 61)
||(x_pointer == 87 && y_pointer == 61)
||(x_pointer == 88 && y_pointer == 61)
||(x_pointer == 89 && y_pointer == 61)
||(x_pointer == 90 && y_pointer == 61)
||(x_pointer == 91 && y_pointer == 61)
||(x_pointer == 155 && y_pointer == 61)
||(x_pointer == 156 && y_pointer == 61)
||(x_pointer == 157 && y_pointer == 61)
||(x_pointer == 2 && y_pointer == 62)
||(x_pointer == 3 && y_pointer == 62)
||(x_pointer == 4 && y_pointer == 62)
||(x_pointer == 56 && y_pointer == 62)
||(x_pointer == 57 && y_pointer == 62)
||(x_pointer == 58 && y_pointer == 62)
||(x_pointer == 59 && y_pointer == 62)
||(x_pointer == 60 && y_pointer == 62)
||(x_pointer == 61 && y_pointer == 62)
||(x_pointer == 62 && y_pointer == 62)
||(x_pointer == 63 && y_pointer == 62)
||(x_pointer == 64 && y_pointer == 62)
||(x_pointer == 65 && y_pointer == 62)
||(x_pointer == 66 && y_pointer == 62)
||(x_pointer == 67 && y_pointer == 62)
||(x_pointer == 68 && y_pointer == 62)
||(x_pointer == 69 && y_pointer == 62)
||(x_pointer == 70 && y_pointer == 62)
||(x_pointer == 71 && y_pointer == 62)
||(x_pointer == 72 && y_pointer == 62)
||(x_pointer == 73 && y_pointer == 62)
||(x_pointer == 74 && y_pointer == 62)
||(x_pointer == 75 && y_pointer == 62)
||(x_pointer == 76 && y_pointer == 62)
||(x_pointer == 77 && y_pointer == 62)
||(x_pointer == 78 && y_pointer == 62)
||(x_pointer == 79 && y_pointer == 62)
||(x_pointer == 80 && y_pointer == 62)
||(x_pointer == 81 && y_pointer == 62)
||(x_pointer == 82 && y_pointer == 62)
||(x_pointer == 83 && y_pointer == 62)
||(x_pointer == 84 && y_pointer == 62)
||(x_pointer == 85 && y_pointer == 62)
||(x_pointer == 86 && y_pointer == 62)
||(x_pointer == 87 && y_pointer == 62)
||(x_pointer == 88 && y_pointer == 62)
||(x_pointer == 89 && y_pointer == 62)
||(x_pointer == 90 && y_pointer == 62)
||(x_pointer == 91 && y_pointer == 62)
||(x_pointer == 92 && y_pointer == 62)
||(x_pointer == 93 && y_pointer == 62)
||(x_pointer == 94 && y_pointer == 62)
||(x_pointer == 95 && y_pointer == 62)
||(x_pointer == 96 && y_pointer == 62)
||(x_pointer == 97 && y_pointer == 62)
||(x_pointer == 98 && y_pointer == 62)
||(x_pointer == 99 && y_pointer == 62)
||(x_pointer == 100 && y_pointer == 62)
||(x_pointer == 101 && y_pointer == 62)
||(x_pointer == 102 && y_pointer == 62)
||(x_pointer == 103 && y_pointer == 62)
||(x_pointer == 104 && y_pointer == 62)
||(x_pointer == 105 && y_pointer == 62)
||(x_pointer == 106 && y_pointer == 62)
||(x_pointer == 155 && y_pointer == 62)
||(x_pointer == 156 && y_pointer == 62)
||(x_pointer == 157 && y_pointer == 62)
||(x_pointer == 2 && y_pointer == 63)
||(x_pointer == 3 && y_pointer == 63)
||(x_pointer == 4 && y_pointer == 63)
||(x_pointer == 56 && y_pointer == 63)
||(x_pointer == 57 && y_pointer == 63)
||(x_pointer == 58 && y_pointer == 63)
||(x_pointer == 59 && y_pointer == 63)
||(x_pointer == 60 && y_pointer == 63)
||(x_pointer == 61 && y_pointer == 63)
||(x_pointer == 62 && y_pointer == 63)
||(x_pointer == 63 && y_pointer == 63)
||(x_pointer == 64 && y_pointer == 63)
||(x_pointer == 65 && y_pointer == 63)
||(x_pointer == 66 && y_pointer == 63)
||(x_pointer == 67 && y_pointer == 63)
||(x_pointer == 68 && y_pointer == 63)
||(x_pointer == 69 && y_pointer == 63)
||(x_pointer == 70 && y_pointer == 63)
||(x_pointer == 71 && y_pointer == 63)
||(x_pointer == 72 && y_pointer == 63)
||(x_pointer == 73 && y_pointer == 63)
||(x_pointer == 74 && y_pointer == 63)
||(x_pointer == 75 && y_pointer == 63)
||(x_pointer == 76 && y_pointer == 63)
||(x_pointer == 77 && y_pointer == 63)
||(x_pointer == 78 && y_pointer == 63)
||(x_pointer == 79 && y_pointer == 63)
||(x_pointer == 80 && y_pointer == 63)
||(x_pointer == 81 && y_pointer == 63)
||(x_pointer == 82 && y_pointer == 63)
||(x_pointer == 83 && y_pointer == 63)
||(x_pointer == 84 && y_pointer == 63)
||(x_pointer == 85 && y_pointer == 63)
||(x_pointer == 86 && y_pointer == 63)
||(x_pointer == 87 && y_pointer == 63)
||(x_pointer == 88 && y_pointer == 63)
||(x_pointer == 89 && y_pointer == 63)
||(x_pointer == 90 && y_pointer == 63)
||(x_pointer == 91 && y_pointer == 63)
||(x_pointer == 92 && y_pointer == 63)
||(x_pointer == 93 && y_pointer == 63)
||(x_pointer == 94 && y_pointer == 63)
||(x_pointer == 95 && y_pointer == 63)
||(x_pointer == 96 && y_pointer == 63)
||(x_pointer == 97 && y_pointer == 63)
||(x_pointer == 98 && y_pointer == 63)
||(x_pointer == 99 && y_pointer == 63)
||(x_pointer == 100 && y_pointer == 63)
||(x_pointer == 101 && y_pointer == 63)
||(x_pointer == 102 && y_pointer == 63)
||(x_pointer == 103 && y_pointer == 63)
||(x_pointer == 104 && y_pointer == 63)
||(x_pointer == 105 && y_pointer == 63)
||(x_pointer == 106 && y_pointer == 63)
||(x_pointer == 155 && y_pointer == 63)
||(x_pointer == 156 && y_pointer == 63)
||(x_pointer == 157 && y_pointer == 63)
||(x_pointer == 2 && y_pointer == 64)
||(x_pointer == 3 && y_pointer == 64)
||(x_pointer == 4 && y_pointer == 64)
||(x_pointer == 56 && y_pointer == 64)
||(x_pointer == 57 && y_pointer == 64)
||(x_pointer == 58 && y_pointer == 64)
||(x_pointer == 59 && y_pointer == 64)
||(x_pointer == 60 && y_pointer == 64)
||(x_pointer == 61 && y_pointer == 64)
||(x_pointer == 62 && y_pointer == 64)
||(x_pointer == 63 && y_pointer == 64)
||(x_pointer == 64 && y_pointer == 64)
||(x_pointer == 65 && y_pointer == 64)
||(x_pointer == 66 && y_pointer == 64)
||(x_pointer == 67 && y_pointer == 64)
||(x_pointer == 68 && y_pointer == 64)
||(x_pointer == 69 && y_pointer == 64)
||(x_pointer == 70 && y_pointer == 64)
||(x_pointer == 71 && y_pointer == 64)
||(x_pointer == 72 && y_pointer == 64)
||(x_pointer == 73 && y_pointer == 64)
||(x_pointer == 74 && y_pointer == 64)
||(x_pointer == 75 && y_pointer == 64)
||(x_pointer == 76 && y_pointer == 64)
||(x_pointer == 77 && y_pointer == 64)
||(x_pointer == 78 && y_pointer == 64)
||(x_pointer == 79 && y_pointer == 64)
||(x_pointer == 80 && y_pointer == 64)
||(x_pointer == 81 && y_pointer == 64)
||(x_pointer == 82 && y_pointer == 64)
||(x_pointer == 83 && y_pointer == 64)
||(x_pointer == 84 && y_pointer == 64)
||(x_pointer == 85 && y_pointer == 64)
||(x_pointer == 86 && y_pointer == 64)
||(x_pointer == 87 && y_pointer == 64)
||(x_pointer == 88 && y_pointer == 64)
||(x_pointer == 89 && y_pointer == 64)
||(x_pointer == 90 && y_pointer == 64)
||(x_pointer == 91 && y_pointer == 64)
||(x_pointer == 92 && y_pointer == 64)
||(x_pointer == 93 && y_pointer == 64)
||(x_pointer == 94 && y_pointer == 64)
||(x_pointer == 95 && y_pointer == 64)
||(x_pointer == 96 && y_pointer == 64)
||(x_pointer == 97 && y_pointer == 64)
||(x_pointer == 98 && y_pointer == 64)
||(x_pointer == 99 && y_pointer == 64)
||(x_pointer == 100 && y_pointer == 64)
||(x_pointer == 101 && y_pointer == 64)
||(x_pointer == 102 && y_pointer == 64)
||(x_pointer == 103 && y_pointer == 64)
||(x_pointer == 104 && y_pointer == 64)
||(x_pointer == 105 && y_pointer == 64)
||(x_pointer == 106 && y_pointer == 64)
||(x_pointer == 155 && y_pointer == 64)
||(x_pointer == 156 && y_pointer == 64)
||(x_pointer == 157 && y_pointer == 64)
||(x_pointer == 2 && y_pointer == 65)
||(x_pointer == 3 && y_pointer == 65)
||(x_pointer == 4 && y_pointer == 65)
||(x_pointer == 56 && y_pointer == 65)
||(x_pointer == 57 && y_pointer == 65)
||(x_pointer == 58 && y_pointer == 65)
||(x_pointer == 59 && y_pointer == 65)
||(x_pointer == 60 && y_pointer == 65)
||(x_pointer == 61 && y_pointer == 65)
||(x_pointer == 62 && y_pointer == 65)
||(x_pointer == 63 && y_pointer == 65)
||(x_pointer == 64 && y_pointer == 65)
||(x_pointer == 65 && y_pointer == 65)
||(x_pointer == 66 && y_pointer == 65)
||(x_pointer == 67 && y_pointer == 65)
||(x_pointer == 68 && y_pointer == 65)
||(x_pointer == 69 && y_pointer == 65)
||(x_pointer == 70 && y_pointer == 65)
||(x_pointer == 71 && y_pointer == 65)
||(x_pointer == 72 && y_pointer == 65)
||(x_pointer == 73 && y_pointer == 65)
||(x_pointer == 74 && y_pointer == 65)
||(x_pointer == 75 && y_pointer == 65)
||(x_pointer == 76 && y_pointer == 65)
||(x_pointer == 77 && y_pointer == 65)
||(x_pointer == 78 && y_pointer == 65)
||(x_pointer == 79 && y_pointer == 65)
||(x_pointer == 80 && y_pointer == 65)
||(x_pointer == 81 && y_pointer == 65)
||(x_pointer == 82 && y_pointer == 65)
||(x_pointer == 83 && y_pointer == 65)
||(x_pointer == 84 && y_pointer == 65)
||(x_pointer == 85 && y_pointer == 65)
||(x_pointer == 86 && y_pointer == 65)
||(x_pointer == 87 && y_pointer == 65)
||(x_pointer == 88 && y_pointer == 65)
||(x_pointer == 89 && y_pointer == 65)
||(x_pointer == 90 && y_pointer == 65)
||(x_pointer == 91 && y_pointer == 65)
||(x_pointer == 92 && y_pointer == 65)
||(x_pointer == 93 && y_pointer == 65)
||(x_pointer == 94 && y_pointer == 65)
||(x_pointer == 95 && y_pointer == 65)
||(x_pointer == 96 && y_pointer == 65)
||(x_pointer == 97 && y_pointer == 65)
||(x_pointer == 98 && y_pointer == 65)
||(x_pointer == 99 && y_pointer == 65)
||(x_pointer == 100 && y_pointer == 65)
||(x_pointer == 101 && y_pointer == 65)
||(x_pointer == 102 && y_pointer == 65)
||(x_pointer == 103 && y_pointer == 65)
||(x_pointer == 104 && y_pointer == 65)
||(x_pointer == 105 && y_pointer == 65)
||(x_pointer == 106 && y_pointer == 65)
||(x_pointer == 155 && y_pointer == 65)
||(x_pointer == 156 && y_pointer == 65)
||(x_pointer == 157 && y_pointer == 65)
||(x_pointer == 2 && y_pointer == 66)
||(x_pointer == 3 && y_pointer == 66)
||(x_pointer == 4 && y_pointer == 66)
||(x_pointer == 56 && y_pointer == 66)
||(x_pointer == 57 && y_pointer == 66)
||(x_pointer == 58 && y_pointer == 66)
||(x_pointer == 59 && y_pointer == 66)
||(x_pointer == 60 && y_pointer == 66)
||(x_pointer == 61 && y_pointer == 66)
||(x_pointer == 62 && y_pointer == 66)
||(x_pointer == 63 && y_pointer == 66)
||(x_pointer == 64 && y_pointer == 66)
||(x_pointer == 65 && y_pointer == 66)
||(x_pointer == 66 && y_pointer == 66)
||(x_pointer == 67 && y_pointer == 66)
||(x_pointer == 68 && y_pointer == 66)
||(x_pointer == 69 && y_pointer == 66)
||(x_pointer == 70 && y_pointer == 66)
||(x_pointer == 71 && y_pointer == 66)
||(x_pointer == 72 && y_pointer == 66)
||(x_pointer == 73 && y_pointer == 66)
||(x_pointer == 74 && y_pointer == 66)
||(x_pointer == 75 && y_pointer == 66)
||(x_pointer == 76 && y_pointer == 66)
||(x_pointer == 77 && y_pointer == 66)
||(x_pointer == 78 && y_pointer == 66)
||(x_pointer == 79 && y_pointer == 66)
||(x_pointer == 80 && y_pointer == 66)
||(x_pointer == 81 && y_pointer == 66)
||(x_pointer == 82 && y_pointer == 66)
||(x_pointer == 83 && y_pointer == 66)
||(x_pointer == 84 && y_pointer == 66)
||(x_pointer == 85 && y_pointer == 66)
||(x_pointer == 86 && y_pointer == 66)
||(x_pointer == 87 && y_pointer == 66)
||(x_pointer == 88 && y_pointer == 66)
||(x_pointer == 89 && y_pointer == 66)
||(x_pointer == 90 && y_pointer == 66)
||(x_pointer == 91 && y_pointer == 66)
||(x_pointer == 92 && y_pointer == 66)
||(x_pointer == 93 && y_pointer == 66)
||(x_pointer == 94 && y_pointer == 66)
||(x_pointer == 95 && y_pointer == 66)
||(x_pointer == 96 && y_pointer == 66)
||(x_pointer == 97 && y_pointer == 66)
||(x_pointer == 98 && y_pointer == 66)
||(x_pointer == 99 && y_pointer == 66)
||(x_pointer == 100 && y_pointer == 66)
||(x_pointer == 101 && y_pointer == 66)
||(x_pointer == 102 && y_pointer == 66)
||(x_pointer == 103 && y_pointer == 66)
||(x_pointer == 104 && y_pointer == 66)
||(x_pointer == 105 && y_pointer == 66)
||(x_pointer == 106 && y_pointer == 66)
||(x_pointer == 155 && y_pointer == 66)
||(x_pointer == 156 && y_pointer == 66)
||(x_pointer == 157 && y_pointer == 66)
||(x_pointer == 2 && y_pointer == 67)
||(x_pointer == 3 && y_pointer == 67)
||(x_pointer == 4 && y_pointer == 67)
||(x_pointer == 56 && y_pointer == 67)
||(x_pointer == 57 && y_pointer == 67)
||(x_pointer == 58 && y_pointer == 67)
||(x_pointer == 59 && y_pointer == 67)
||(x_pointer == 60 && y_pointer == 67)
||(x_pointer == 61 && y_pointer == 67)
||(x_pointer == 62 && y_pointer == 67)
||(x_pointer == 63 && y_pointer == 67)
||(x_pointer == 64 && y_pointer == 67)
||(x_pointer == 65 && y_pointer == 67)
||(x_pointer == 66 && y_pointer == 67)
||(x_pointer == 67 && y_pointer == 67)
||(x_pointer == 68 && y_pointer == 67)
||(x_pointer == 69 && y_pointer == 67)
||(x_pointer == 70 && y_pointer == 67)
||(x_pointer == 71 && y_pointer == 67)
||(x_pointer == 72 && y_pointer == 67)
||(x_pointer == 73 && y_pointer == 67)
||(x_pointer == 74 && y_pointer == 67)
||(x_pointer == 75 && y_pointer == 67)
||(x_pointer == 76 && y_pointer == 67)
||(x_pointer == 77 && y_pointer == 67)
||(x_pointer == 78 && y_pointer == 67)
||(x_pointer == 79 && y_pointer == 67)
||(x_pointer == 80 && y_pointer == 67)
||(x_pointer == 81 && y_pointer == 67)
||(x_pointer == 82 && y_pointer == 67)
||(x_pointer == 83 && y_pointer == 67)
||(x_pointer == 84 && y_pointer == 67)
||(x_pointer == 85 && y_pointer == 67)
||(x_pointer == 86 && y_pointer == 67)
||(x_pointer == 87 && y_pointer == 67)
||(x_pointer == 88 && y_pointer == 67)
||(x_pointer == 89 && y_pointer == 67)
||(x_pointer == 90 && y_pointer == 67)
||(x_pointer == 91 && y_pointer == 67)
||(x_pointer == 92 && y_pointer == 67)
||(x_pointer == 93 && y_pointer == 67)
||(x_pointer == 94 && y_pointer == 67)
||(x_pointer == 95 && y_pointer == 67)
||(x_pointer == 96 && y_pointer == 67)
||(x_pointer == 97 && y_pointer == 67)
||(x_pointer == 98 && y_pointer == 67)
||(x_pointer == 99 && y_pointer == 67)
||(x_pointer == 100 && y_pointer == 67)
||(x_pointer == 101 && y_pointer == 67)
||(x_pointer == 102 && y_pointer == 67)
||(x_pointer == 103 && y_pointer == 67)
||(x_pointer == 104 && y_pointer == 67)
||(x_pointer == 105 && y_pointer == 67)
||(x_pointer == 106 && y_pointer == 67)
||(x_pointer == 155 && y_pointer == 67)
||(x_pointer == 156 && y_pointer == 67)
||(x_pointer == 157 && y_pointer == 67)
||(x_pointer == 2 && y_pointer == 68)
||(x_pointer == 3 && y_pointer == 68)
||(x_pointer == 4 && y_pointer == 68)
||(x_pointer == 56 && y_pointer == 68)
||(x_pointer == 57 && y_pointer == 68)
||(x_pointer == 58 && y_pointer == 68)
||(x_pointer == 59 && y_pointer == 68)
||(x_pointer == 60 && y_pointer == 68)
||(x_pointer == 61 && y_pointer == 68)
||(x_pointer == 62 && y_pointer == 68)
||(x_pointer == 63 && y_pointer == 68)
||(x_pointer == 64 && y_pointer == 68)
||(x_pointer == 65 && y_pointer == 68)
||(x_pointer == 66 && y_pointer == 68)
||(x_pointer == 67 && y_pointer == 68)
||(x_pointer == 68 && y_pointer == 68)
||(x_pointer == 69 && y_pointer == 68)
||(x_pointer == 70 && y_pointer == 68)
||(x_pointer == 71 && y_pointer == 68)
||(x_pointer == 72 && y_pointer == 68)
||(x_pointer == 73 && y_pointer == 68)
||(x_pointer == 74 && y_pointer == 68)
||(x_pointer == 75 && y_pointer == 68)
||(x_pointer == 76 && y_pointer == 68)
||(x_pointer == 77 && y_pointer == 68)
||(x_pointer == 78 && y_pointer == 68)
||(x_pointer == 79 && y_pointer == 68)
||(x_pointer == 80 && y_pointer == 68)
||(x_pointer == 81 && y_pointer == 68)
||(x_pointer == 82 && y_pointer == 68)
||(x_pointer == 83 && y_pointer == 68)
||(x_pointer == 84 && y_pointer == 68)
||(x_pointer == 85 && y_pointer == 68)
||(x_pointer == 86 && y_pointer == 68)
||(x_pointer == 87 && y_pointer == 68)
||(x_pointer == 88 && y_pointer == 68)
||(x_pointer == 89 && y_pointer == 68)
||(x_pointer == 90 && y_pointer == 68)
||(x_pointer == 91 && y_pointer == 68)
||(x_pointer == 92 && y_pointer == 68)
||(x_pointer == 93 && y_pointer == 68)
||(x_pointer == 94 && y_pointer == 68)
||(x_pointer == 95 && y_pointer == 68)
||(x_pointer == 96 && y_pointer == 68)
||(x_pointer == 97 && y_pointer == 68)
||(x_pointer == 98 && y_pointer == 68)
||(x_pointer == 99 && y_pointer == 68)
||(x_pointer == 100 && y_pointer == 68)
||(x_pointer == 101 && y_pointer == 68)
||(x_pointer == 102 && y_pointer == 68)
||(x_pointer == 103 && y_pointer == 68)
||(x_pointer == 104 && y_pointer == 68)
||(x_pointer == 105 && y_pointer == 68)
||(x_pointer == 106 && y_pointer == 68)
||(x_pointer == 155 && y_pointer == 68)
||(x_pointer == 156 && y_pointer == 68)
||(x_pointer == 157 && y_pointer == 68)
||(x_pointer == 2 && y_pointer == 69)
||(x_pointer == 3 && y_pointer == 69)
||(x_pointer == 4 && y_pointer == 69)
||(x_pointer == 56 && y_pointer == 69)
||(x_pointer == 57 && y_pointer == 69)
||(x_pointer == 58 && y_pointer == 69)
||(x_pointer == 59 && y_pointer == 69)
||(x_pointer == 60 && y_pointer == 69)
||(x_pointer == 61 && y_pointer == 69)
||(x_pointer == 62 && y_pointer == 69)
||(x_pointer == 63 && y_pointer == 69)
||(x_pointer == 64 && y_pointer == 69)
||(x_pointer == 65 && y_pointer == 69)
||(x_pointer == 66 && y_pointer == 69)
||(x_pointer == 67 && y_pointer == 69)
||(x_pointer == 68 && y_pointer == 69)
||(x_pointer == 69 && y_pointer == 69)
||(x_pointer == 70 && y_pointer == 69)
||(x_pointer == 71 && y_pointer == 69)
||(x_pointer == 72 && y_pointer == 69)
||(x_pointer == 73 && y_pointer == 69)
||(x_pointer == 74 && y_pointer == 69)
||(x_pointer == 75 && y_pointer == 69)
||(x_pointer == 76 && y_pointer == 69)
||(x_pointer == 77 && y_pointer == 69)
||(x_pointer == 78 && y_pointer == 69)
||(x_pointer == 79 && y_pointer == 69)
||(x_pointer == 80 && y_pointer == 69)
||(x_pointer == 81 && y_pointer == 69)
||(x_pointer == 82 && y_pointer == 69)
||(x_pointer == 83 && y_pointer == 69)
||(x_pointer == 84 && y_pointer == 69)
||(x_pointer == 85 && y_pointer == 69)
||(x_pointer == 86 && y_pointer == 69)
||(x_pointer == 87 && y_pointer == 69)
||(x_pointer == 88 && y_pointer == 69)
||(x_pointer == 89 && y_pointer == 69)
||(x_pointer == 90 && y_pointer == 69)
||(x_pointer == 91 && y_pointer == 69)
||(x_pointer == 92 && y_pointer == 69)
||(x_pointer == 93 && y_pointer == 69)
||(x_pointer == 94 && y_pointer == 69)
||(x_pointer == 95 && y_pointer == 69)
||(x_pointer == 96 && y_pointer == 69)
||(x_pointer == 97 && y_pointer == 69)
||(x_pointer == 98 && y_pointer == 69)
||(x_pointer == 99 && y_pointer == 69)
||(x_pointer == 100 && y_pointer == 69)
||(x_pointer == 101 && y_pointer == 69)
||(x_pointer == 102 && y_pointer == 69)
||(x_pointer == 103 && y_pointer == 69)
||(x_pointer == 104 && y_pointer == 69)
||(x_pointer == 105 && y_pointer == 69)
||(x_pointer == 106 && y_pointer == 69)
||(x_pointer == 155 && y_pointer == 69)
||(x_pointer == 156 && y_pointer == 69)
||(x_pointer == 157 && y_pointer == 69)
||(x_pointer == 2 && y_pointer == 70)
||(x_pointer == 3 && y_pointer == 70)
||(x_pointer == 4 && y_pointer == 70)
||(x_pointer == 56 && y_pointer == 70)
||(x_pointer == 57 && y_pointer == 70)
||(x_pointer == 58 && y_pointer == 70)
||(x_pointer == 59 && y_pointer == 70)
||(x_pointer == 60 && y_pointer == 70)
||(x_pointer == 61 && y_pointer == 70)
||(x_pointer == 62 && y_pointer == 70)
||(x_pointer == 63 && y_pointer == 70)
||(x_pointer == 64 && y_pointer == 70)
||(x_pointer == 65 && y_pointer == 70)
||(x_pointer == 66 && y_pointer == 70)
||(x_pointer == 67 && y_pointer == 70)
||(x_pointer == 68 && y_pointer == 70)
||(x_pointer == 69 && y_pointer == 70)
||(x_pointer == 70 && y_pointer == 70)
||(x_pointer == 71 && y_pointer == 70)
||(x_pointer == 72 && y_pointer == 70)
||(x_pointer == 73 && y_pointer == 70)
||(x_pointer == 74 && y_pointer == 70)
||(x_pointer == 75 && y_pointer == 70)
||(x_pointer == 76 && y_pointer == 70)
||(x_pointer == 77 && y_pointer == 70)
||(x_pointer == 78 && y_pointer == 70)
||(x_pointer == 79 && y_pointer == 70)
||(x_pointer == 80 && y_pointer == 70)
||(x_pointer == 81 && y_pointer == 70)
||(x_pointer == 82 && y_pointer == 70)
||(x_pointer == 83 && y_pointer == 70)
||(x_pointer == 84 && y_pointer == 70)
||(x_pointer == 85 && y_pointer == 70)
||(x_pointer == 86 && y_pointer == 70)
||(x_pointer == 87 && y_pointer == 70)
||(x_pointer == 88 && y_pointer == 70)
||(x_pointer == 89 && y_pointer == 70)
||(x_pointer == 90 && y_pointer == 70)
||(x_pointer == 91 && y_pointer == 70)
||(x_pointer == 92 && y_pointer == 70)
||(x_pointer == 93 && y_pointer == 70)
||(x_pointer == 94 && y_pointer == 70)
||(x_pointer == 95 && y_pointer == 70)
||(x_pointer == 96 && y_pointer == 70)
||(x_pointer == 97 && y_pointer == 70)
||(x_pointer == 98 && y_pointer == 70)
||(x_pointer == 99 && y_pointer == 70)
||(x_pointer == 100 && y_pointer == 70)
||(x_pointer == 101 && y_pointer == 70)
||(x_pointer == 102 && y_pointer == 70)
||(x_pointer == 103 && y_pointer == 70)
||(x_pointer == 104 && y_pointer == 70)
||(x_pointer == 105 && y_pointer == 70)
||(x_pointer == 106 && y_pointer == 70)
||(x_pointer == 155 && y_pointer == 70)
||(x_pointer == 156 && y_pointer == 70)
||(x_pointer == 157 && y_pointer == 70)
||(x_pointer == 2 && y_pointer == 71)
||(x_pointer == 3 && y_pointer == 71)
||(x_pointer == 4 && y_pointer == 71)
||(x_pointer == 56 && y_pointer == 71)
||(x_pointer == 57 && y_pointer == 71)
||(x_pointer == 58 && y_pointer == 71)
||(x_pointer == 59 && y_pointer == 71)
||(x_pointer == 60 && y_pointer == 71)
||(x_pointer == 61 && y_pointer == 71)
||(x_pointer == 62 && y_pointer == 71)
||(x_pointer == 63 && y_pointer == 71)
||(x_pointer == 64 && y_pointer == 71)
||(x_pointer == 65 && y_pointer == 71)
||(x_pointer == 66 && y_pointer == 71)
||(x_pointer == 67 && y_pointer == 71)
||(x_pointer == 68 && y_pointer == 71)
||(x_pointer == 69 && y_pointer == 71)
||(x_pointer == 70 && y_pointer == 71)
||(x_pointer == 71 && y_pointer == 71)
||(x_pointer == 72 && y_pointer == 71)
||(x_pointer == 73 && y_pointer == 71)
||(x_pointer == 74 && y_pointer == 71)
||(x_pointer == 75 && y_pointer == 71)
||(x_pointer == 76 && y_pointer == 71)
||(x_pointer == 77 && y_pointer == 71)
||(x_pointer == 78 && y_pointer == 71)
||(x_pointer == 79 && y_pointer == 71)
||(x_pointer == 80 && y_pointer == 71)
||(x_pointer == 81 && y_pointer == 71)
||(x_pointer == 82 && y_pointer == 71)
||(x_pointer == 83 && y_pointer == 71)
||(x_pointer == 84 && y_pointer == 71)
||(x_pointer == 85 && y_pointer == 71)
||(x_pointer == 86 && y_pointer == 71)
||(x_pointer == 87 && y_pointer == 71)
||(x_pointer == 88 && y_pointer == 71)
||(x_pointer == 89 && y_pointer == 71)
||(x_pointer == 90 && y_pointer == 71)
||(x_pointer == 91 && y_pointer == 71)
||(x_pointer == 92 && y_pointer == 71)
||(x_pointer == 93 && y_pointer == 71)
||(x_pointer == 94 && y_pointer == 71)
||(x_pointer == 95 && y_pointer == 71)
||(x_pointer == 96 && y_pointer == 71)
||(x_pointer == 97 && y_pointer == 71)
||(x_pointer == 98 && y_pointer == 71)
||(x_pointer == 99 && y_pointer == 71)
||(x_pointer == 100 && y_pointer == 71)
||(x_pointer == 101 && y_pointer == 71)
||(x_pointer == 102 && y_pointer == 71)
||(x_pointer == 103 && y_pointer == 71)
||(x_pointer == 104 && y_pointer == 71)
||(x_pointer == 105 && y_pointer == 71)
||(x_pointer == 106 && y_pointer == 71)
||(x_pointer == 155 && y_pointer == 71)
||(x_pointer == 156 && y_pointer == 71)
||(x_pointer == 157 && y_pointer == 71)
||(x_pointer == 2 && y_pointer == 72)
||(x_pointer == 3 && y_pointer == 72)
||(x_pointer == 4 && y_pointer == 72)
||(x_pointer == 56 && y_pointer == 72)
||(x_pointer == 57 && y_pointer == 72)
||(x_pointer == 58 && y_pointer == 72)
||(x_pointer == 59 && y_pointer == 72)
||(x_pointer == 60 && y_pointer == 72)
||(x_pointer == 61 && y_pointer == 72)
||(x_pointer == 62 && y_pointer == 72)
||(x_pointer == 63 && y_pointer == 72)
||(x_pointer == 64 && y_pointer == 72)
||(x_pointer == 65 && y_pointer == 72)
||(x_pointer == 66 && y_pointer == 72)
||(x_pointer == 67 && y_pointer == 72)
||(x_pointer == 68 && y_pointer == 72)
||(x_pointer == 69 && y_pointer == 72)
||(x_pointer == 70 && y_pointer == 72)
||(x_pointer == 71 && y_pointer == 72)
||(x_pointer == 72 && y_pointer == 72)
||(x_pointer == 73 && y_pointer == 72)
||(x_pointer == 74 && y_pointer == 72)
||(x_pointer == 75 && y_pointer == 72)
||(x_pointer == 76 && y_pointer == 72)
||(x_pointer == 77 && y_pointer == 72)
||(x_pointer == 78 && y_pointer == 72)
||(x_pointer == 79 && y_pointer == 72)
||(x_pointer == 80 && y_pointer == 72)
||(x_pointer == 81 && y_pointer == 72)
||(x_pointer == 82 && y_pointer == 72)
||(x_pointer == 83 && y_pointer == 72)
||(x_pointer == 84 && y_pointer == 72)
||(x_pointer == 85 && y_pointer == 72)
||(x_pointer == 86 && y_pointer == 72)
||(x_pointer == 87 && y_pointer == 72)
||(x_pointer == 88 && y_pointer == 72)
||(x_pointer == 89 && y_pointer == 72)
||(x_pointer == 90 && y_pointer == 72)
||(x_pointer == 91 && y_pointer == 72)
||(x_pointer == 92 && y_pointer == 72)
||(x_pointer == 93 && y_pointer == 72)
||(x_pointer == 94 && y_pointer == 72)
||(x_pointer == 95 && y_pointer == 72)
||(x_pointer == 96 && y_pointer == 72)
||(x_pointer == 97 && y_pointer == 72)
||(x_pointer == 98 && y_pointer == 72)
||(x_pointer == 99 && y_pointer == 72)
||(x_pointer == 100 && y_pointer == 72)
||(x_pointer == 101 && y_pointer == 72)
||(x_pointer == 102 && y_pointer == 72)
||(x_pointer == 103 && y_pointer == 72)
||(x_pointer == 104 && y_pointer == 72)
||(x_pointer == 105 && y_pointer == 72)
||(x_pointer == 106 && y_pointer == 72)
||(x_pointer == 155 && y_pointer == 72)
||(x_pointer == 156 && y_pointer == 72)
||(x_pointer == 157 && y_pointer == 72)
||(x_pointer == 2 && y_pointer == 73)
||(x_pointer == 3 && y_pointer == 73)
||(x_pointer == 4 && y_pointer == 73)
||(x_pointer == 56 && y_pointer == 73)
||(x_pointer == 57 && y_pointer == 73)
||(x_pointer == 58 && y_pointer == 73)
||(x_pointer == 59 && y_pointer == 73)
||(x_pointer == 60 && y_pointer == 73)
||(x_pointer == 61 && y_pointer == 73)
||(x_pointer == 62 && y_pointer == 73)
||(x_pointer == 63 && y_pointer == 73)
||(x_pointer == 64 && y_pointer == 73)
||(x_pointer == 65 && y_pointer == 73)
||(x_pointer == 66 && y_pointer == 73)
||(x_pointer == 67 && y_pointer == 73)
||(x_pointer == 68 && y_pointer == 73)
||(x_pointer == 69 && y_pointer == 73)
||(x_pointer == 70 && y_pointer == 73)
||(x_pointer == 71 && y_pointer == 73)
||(x_pointer == 72 && y_pointer == 73)
||(x_pointer == 73 && y_pointer == 73)
||(x_pointer == 74 && y_pointer == 73)
||(x_pointer == 75 && y_pointer == 73)
||(x_pointer == 76 && y_pointer == 73)
||(x_pointer == 77 && y_pointer == 73)
||(x_pointer == 78 && y_pointer == 73)
||(x_pointer == 79 && y_pointer == 73)
||(x_pointer == 80 && y_pointer == 73)
||(x_pointer == 81 && y_pointer == 73)
||(x_pointer == 82 && y_pointer == 73)
||(x_pointer == 83 && y_pointer == 73)
||(x_pointer == 84 && y_pointer == 73)
||(x_pointer == 85 && y_pointer == 73)
||(x_pointer == 86 && y_pointer == 73)
||(x_pointer == 87 && y_pointer == 73)
||(x_pointer == 88 && y_pointer == 73)
||(x_pointer == 89 && y_pointer == 73)
||(x_pointer == 90 && y_pointer == 73)
||(x_pointer == 91 && y_pointer == 73)
||(x_pointer == 92 && y_pointer == 73)
||(x_pointer == 93 && y_pointer == 73)
||(x_pointer == 94 && y_pointer == 73)
||(x_pointer == 95 && y_pointer == 73)
||(x_pointer == 96 && y_pointer == 73)
||(x_pointer == 97 && y_pointer == 73)
||(x_pointer == 98 && y_pointer == 73)
||(x_pointer == 99 && y_pointer == 73)
||(x_pointer == 100 && y_pointer == 73)
||(x_pointer == 101 && y_pointer == 73)
||(x_pointer == 102 && y_pointer == 73)
||(x_pointer == 103 && y_pointer == 73)
||(x_pointer == 104 && y_pointer == 73)
||(x_pointer == 105 && y_pointer == 73)
||(x_pointer == 106 && y_pointer == 73)
||(x_pointer == 155 && y_pointer == 73)
||(x_pointer == 156 && y_pointer == 73)
||(x_pointer == 157 && y_pointer == 73)
||(x_pointer == 2 && y_pointer == 74)
||(x_pointer == 3 && y_pointer == 74)
||(x_pointer == 4 && y_pointer == 74)
||(x_pointer == 56 && y_pointer == 74)
||(x_pointer == 57 && y_pointer == 74)
||(x_pointer == 58 && y_pointer == 74)
||(x_pointer == 59 && y_pointer == 74)
||(x_pointer == 60 && y_pointer == 74)
||(x_pointer == 61 && y_pointer == 74)
||(x_pointer == 62 && y_pointer == 74)
||(x_pointer == 63 && y_pointer == 74)
||(x_pointer == 64 && y_pointer == 74)
||(x_pointer == 65 && y_pointer == 74)
||(x_pointer == 66 && y_pointer == 74)
||(x_pointer == 67 && y_pointer == 74)
||(x_pointer == 68 && y_pointer == 74)
||(x_pointer == 69 && y_pointer == 74)
||(x_pointer == 70 && y_pointer == 74)
||(x_pointer == 71 && y_pointer == 74)
||(x_pointer == 72 && y_pointer == 74)
||(x_pointer == 73 && y_pointer == 74)
||(x_pointer == 74 && y_pointer == 74)
||(x_pointer == 75 && y_pointer == 74)
||(x_pointer == 76 && y_pointer == 74)
||(x_pointer == 77 && y_pointer == 74)
||(x_pointer == 78 && y_pointer == 74)
||(x_pointer == 79 && y_pointer == 74)
||(x_pointer == 80 && y_pointer == 74)
||(x_pointer == 81 && y_pointer == 74)
||(x_pointer == 82 && y_pointer == 74)
||(x_pointer == 83 && y_pointer == 74)
||(x_pointer == 84 && y_pointer == 74)
||(x_pointer == 85 && y_pointer == 74)
||(x_pointer == 86 && y_pointer == 74)
||(x_pointer == 87 && y_pointer == 74)
||(x_pointer == 88 && y_pointer == 74)
||(x_pointer == 89 && y_pointer == 74)
||(x_pointer == 90 && y_pointer == 74)
||(x_pointer == 91 && y_pointer == 74)
||(x_pointer == 92 && y_pointer == 74)
||(x_pointer == 93 && y_pointer == 74)
||(x_pointer == 94 && y_pointer == 74)
||(x_pointer == 95 && y_pointer == 74)
||(x_pointer == 96 && y_pointer == 74)
||(x_pointer == 97 && y_pointer == 74)
||(x_pointer == 98 && y_pointer == 74)
||(x_pointer == 99 && y_pointer == 74)
||(x_pointer == 100 && y_pointer == 74)
||(x_pointer == 101 && y_pointer == 74)
||(x_pointer == 102 && y_pointer == 74)
||(x_pointer == 103 && y_pointer == 74)
||(x_pointer == 104 && y_pointer == 74)
||(x_pointer == 105 && y_pointer == 74)
||(x_pointer == 106 && y_pointer == 74)
||(x_pointer == 155 && y_pointer == 74)
||(x_pointer == 156 && y_pointer == 74)
||(x_pointer == 157 && y_pointer == 74)
||(x_pointer == 2 && y_pointer == 75)
||(x_pointer == 3 && y_pointer == 75)
||(x_pointer == 4 && y_pointer == 75)
||(x_pointer == 56 && y_pointer == 75)
||(x_pointer == 57 && y_pointer == 75)
||(x_pointer == 58 && y_pointer == 75)
||(x_pointer == 59 && y_pointer == 75)
||(x_pointer == 60 && y_pointer == 75)
||(x_pointer == 61 && y_pointer == 75)
||(x_pointer == 62 && y_pointer == 75)
||(x_pointer == 63 && y_pointer == 75)
||(x_pointer == 64 && y_pointer == 75)
||(x_pointer == 65 && y_pointer == 75)
||(x_pointer == 66 && y_pointer == 75)
||(x_pointer == 67 && y_pointer == 75)
||(x_pointer == 68 && y_pointer == 75)
||(x_pointer == 69 && y_pointer == 75)
||(x_pointer == 70 && y_pointer == 75)
||(x_pointer == 71 && y_pointer == 75)
||(x_pointer == 72 && y_pointer == 75)
||(x_pointer == 73 && y_pointer == 75)
||(x_pointer == 74 && y_pointer == 75)
||(x_pointer == 75 && y_pointer == 75)
||(x_pointer == 76 && y_pointer == 75)
||(x_pointer == 77 && y_pointer == 75)
||(x_pointer == 78 && y_pointer == 75)
||(x_pointer == 79 && y_pointer == 75)
||(x_pointer == 80 && y_pointer == 75)
||(x_pointer == 81 && y_pointer == 75)
||(x_pointer == 82 && y_pointer == 75)
||(x_pointer == 83 && y_pointer == 75)
||(x_pointer == 84 && y_pointer == 75)
||(x_pointer == 85 && y_pointer == 75)
||(x_pointer == 86 && y_pointer == 75)
||(x_pointer == 87 && y_pointer == 75)
||(x_pointer == 88 && y_pointer == 75)
||(x_pointer == 89 && y_pointer == 75)
||(x_pointer == 90 && y_pointer == 75)
||(x_pointer == 91 && y_pointer == 75)
||(x_pointer == 92 && y_pointer == 75)
||(x_pointer == 93 && y_pointer == 75)
||(x_pointer == 94 && y_pointer == 75)
||(x_pointer == 95 && y_pointer == 75)
||(x_pointer == 96 && y_pointer == 75)
||(x_pointer == 97 && y_pointer == 75)
||(x_pointer == 98 && y_pointer == 75)
||(x_pointer == 99 && y_pointer == 75)
||(x_pointer == 100 && y_pointer == 75)
||(x_pointer == 101 && y_pointer == 75)
||(x_pointer == 102 && y_pointer == 75)
||(x_pointer == 103 && y_pointer == 75)
||(x_pointer == 104 && y_pointer == 75)
||(x_pointer == 105 && y_pointer == 75)
||(x_pointer == 106 && y_pointer == 75)
||(x_pointer == 155 && y_pointer == 75)
||(x_pointer == 156 && y_pointer == 75)
||(x_pointer == 157 && y_pointer == 75)
||(x_pointer == 2 && y_pointer == 76)
||(x_pointer == 3 && y_pointer == 76)
||(x_pointer == 4 && y_pointer == 76)
||(x_pointer == 56 && y_pointer == 76)
||(x_pointer == 57 && y_pointer == 76)
||(x_pointer == 58 && y_pointer == 76)
||(x_pointer == 59 && y_pointer == 76)
||(x_pointer == 60 && y_pointer == 76)
||(x_pointer == 61 && y_pointer == 76)
||(x_pointer == 62 && y_pointer == 76)
||(x_pointer == 63 && y_pointer == 76)
||(x_pointer == 64 && y_pointer == 76)
||(x_pointer == 65 && y_pointer == 76)
||(x_pointer == 66 && y_pointer == 76)
||(x_pointer == 67 && y_pointer == 76)
||(x_pointer == 68 && y_pointer == 76)
||(x_pointer == 69 && y_pointer == 76)
||(x_pointer == 70 && y_pointer == 76)
||(x_pointer == 71 && y_pointer == 76)
||(x_pointer == 72 && y_pointer == 76)
||(x_pointer == 73 && y_pointer == 76)
||(x_pointer == 74 && y_pointer == 76)
||(x_pointer == 75 && y_pointer == 76)
||(x_pointer == 76 && y_pointer == 76)
||(x_pointer == 77 && y_pointer == 76)
||(x_pointer == 78 && y_pointer == 76)
||(x_pointer == 79 && y_pointer == 76)
||(x_pointer == 80 && y_pointer == 76)
||(x_pointer == 81 && y_pointer == 76)
||(x_pointer == 82 && y_pointer == 76)
||(x_pointer == 83 && y_pointer == 76)
||(x_pointer == 84 && y_pointer == 76)
||(x_pointer == 85 && y_pointer == 76)
||(x_pointer == 86 && y_pointer == 76)
||(x_pointer == 87 && y_pointer == 76)
||(x_pointer == 88 && y_pointer == 76)
||(x_pointer == 89 && y_pointer == 76)
||(x_pointer == 90 && y_pointer == 76)
||(x_pointer == 91 && y_pointer == 76)
||(x_pointer == 92 && y_pointer == 76)
||(x_pointer == 93 && y_pointer == 76)
||(x_pointer == 94 && y_pointer == 76)
||(x_pointer == 95 && y_pointer == 76)
||(x_pointer == 96 && y_pointer == 76)
||(x_pointer == 97 && y_pointer == 76)
||(x_pointer == 98 && y_pointer == 76)
||(x_pointer == 99 && y_pointer == 76)
||(x_pointer == 100 && y_pointer == 76)
||(x_pointer == 101 && y_pointer == 76)
||(x_pointer == 102 && y_pointer == 76)
||(x_pointer == 103 && y_pointer == 76)
||(x_pointer == 104 && y_pointer == 76)
||(x_pointer == 105 && y_pointer == 76)
||(x_pointer == 106 && y_pointer == 76)
||(x_pointer == 155 && y_pointer == 76)
||(x_pointer == 156 && y_pointer == 76)
||(x_pointer == 157 && y_pointer == 76)
||(x_pointer == 2 && y_pointer == 77)
||(x_pointer == 3 && y_pointer == 77)
||(x_pointer == 4 && y_pointer == 77)
||(x_pointer == 56 && y_pointer == 77)
||(x_pointer == 57 && y_pointer == 77)
||(x_pointer == 58 && y_pointer == 77)
||(x_pointer == 59 && y_pointer == 77)
||(x_pointer == 60 && y_pointer == 77)
||(x_pointer == 61 && y_pointer == 77)
||(x_pointer == 62 && y_pointer == 77)
||(x_pointer == 63 && y_pointer == 77)
||(x_pointer == 64 && y_pointer == 77)
||(x_pointer == 65 && y_pointer == 77)
||(x_pointer == 66 && y_pointer == 77)
||(x_pointer == 67 && y_pointer == 77)
||(x_pointer == 68 && y_pointer == 77)
||(x_pointer == 69 && y_pointer == 77)
||(x_pointer == 70 && y_pointer == 77)
||(x_pointer == 71 && y_pointer == 77)
||(x_pointer == 72 && y_pointer == 77)
||(x_pointer == 73 && y_pointer == 77)
||(x_pointer == 74 && y_pointer == 77)
||(x_pointer == 75 && y_pointer == 77)
||(x_pointer == 76 && y_pointer == 77)
||(x_pointer == 77 && y_pointer == 77)
||(x_pointer == 78 && y_pointer == 77)
||(x_pointer == 79 && y_pointer == 77)
||(x_pointer == 80 && y_pointer == 77)
||(x_pointer == 81 && y_pointer == 77)
||(x_pointer == 82 && y_pointer == 77)
||(x_pointer == 83 && y_pointer == 77)
||(x_pointer == 84 && y_pointer == 77)
||(x_pointer == 85 && y_pointer == 77)
||(x_pointer == 86 && y_pointer == 77)
||(x_pointer == 87 && y_pointer == 77)
||(x_pointer == 88 && y_pointer == 77)
||(x_pointer == 89 && y_pointer == 77)
||(x_pointer == 90 && y_pointer == 77)
||(x_pointer == 91 && y_pointer == 77)
||(x_pointer == 92 && y_pointer == 77)
||(x_pointer == 93 && y_pointer == 77)
||(x_pointer == 94 && y_pointer == 77)
||(x_pointer == 95 && y_pointer == 77)
||(x_pointer == 96 && y_pointer == 77)
||(x_pointer == 97 && y_pointer == 77)
||(x_pointer == 98 && y_pointer == 77)
||(x_pointer == 99 && y_pointer == 77)
||(x_pointer == 100 && y_pointer == 77)
||(x_pointer == 101 && y_pointer == 77)
||(x_pointer == 102 && y_pointer == 77)
||(x_pointer == 103 && y_pointer == 77)
||(x_pointer == 104 && y_pointer == 77)
||(x_pointer == 105 && y_pointer == 77)
||(x_pointer == 106 && y_pointer == 77)
||(x_pointer == 155 && y_pointer == 77)
||(x_pointer == 156 && y_pointer == 77)
||(x_pointer == 157 && y_pointer == 77)
||(x_pointer == 2 && y_pointer == 78)
||(x_pointer == 3 && y_pointer == 78)
||(x_pointer == 4 && y_pointer == 78)
||(x_pointer == 56 && y_pointer == 78)
||(x_pointer == 57 && y_pointer == 78)
||(x_pointer == 58 && y_pointer == 78)
||(x_pointer == 59 && y_pointer == 78)
||(x_pointer == 60 && y_pointer == 78)
||(x_pointer == 61 && y_pointer == 78)
||(x_pointer == 62 && y_pointer == 78)
||(x_pointer == 63 && y_pointer == 78)
||(x_pointer == 64 && y_pointer == 78)
||(x_pointer == 65 && y_pointer == 78)
||(x_pointer == 66 && y_pointer == 78)
||(x_pointer == 67 && y_pointer == 78)
||(x_pointer == 68 && y_pointer == 78)
||(x_pointer == 69 && y_pointer == 78)
||(x_pointer == 70 && y_pointer == 78)
||(x_pointer == 71 && y_pointer == 78)
||(x_pointer == 72 && y_pointer == 78)
||(x_pointer == 73 && y_pointer == 78)
||(x_pointer == 74 && y_pointer == 78)
||(x_pointer == 75 && y_pointer == 78)
||(x_pointer == 76 && y_pointer == 78)
||(x_pointer == 77 && y_pointer == 78)
||(x_pointer == 78 && y_pointer == 78)
||(x_pointer == 79 && y_pointer == 78)
||(x_pointer == 80 && y_pointer == 78)
||(x_pointer == 81 && y_pointer == 78)
||(x_pointer == 82 && y_pointer == 78)
||(x_pointer == 83 && y_pointer == 78)
||(x_pointer == 84 && y_pointer == 78)
||(x_pointer == 85 && y_pointer == 78)
||(x_pointer == 86 && y_pointer == 78)
||(x_pointer == 87 && y_pointer == 78)
||(x_pointer == 88 && y_pointer == 78)
||(x_pointer == 89 && y_pointer == 78)
||(x_pointer == 90 && y_pointer == 78)
||(x_pointer == 91 && y_pointer == 78)
||(x_pointer == 92 && y_pointer == 78)
||(x_pointer == 93 && y_pointer == 78)
||(x_pointer == 94 && y_pointer == 78)
||(x_pointer == 95 && y_pointer == 78)
||(x_pointer == 96 && y_pointer == 78)
||(x_pointer == 97 && y_pointer == 78)
||(x_pointer == 98 && y_pointer == 78)
||(x_pointer == 99 && y_pointer == 78)
||(x_pointer == 100 && y_pointer == 78)
||(x_pointer == 101 && y_pointer == 78)
||(x_pointer == 102 && y_pointer == 78)
||(x_pointer == 103 && y_pointer == 78)
||(x_pointer == 104 && y_pointer == 78)
||(x_pointer == 105 && y_pointer == 78)
||(x_pointer == 106 && y_pointer == 78)
||(x_pointer == 155 && y_pointer == 78)
||(x_pointer == 156 && y_pointer == 78)
||(x_pointer == 157 && y_pointer == 78)
||(x_pointer == 2 && y_pointer == 79)
||(x_pointer == 3 && y_pointer == 79)
||(x_pointer == 4 && y_pointer == 79)
||(x_pointer == 56 && y_pointer == 79)
||(x_pointer == 57 && y_pointer == 79)
||(x_pointer == 58 && y_pointer == 79)
||(x_pointer == 59 && y_pointer == 79)
||(x_pointer == 60 && y_pointer == 79)
||(x_pointer == 61 && y_pointer == 79)
||(x_pointer == 62 && y_pointer == 79)
||(x_pointer == 63 && y_pointer == 79)
||(x_pointer == 64 && y_pointer == 79)
||(x_pointer == 65 && y_pointer == 79)
||(x_pointer == 66 && y_pointer == 79)
||(x_pointer == 67 && y_pointer == 79)
||(x_pointer == 68 && y_pointer == 79)
||(x_pointer == 69 && y_pointer == 79)
||(x_pointer == 70 && y_pointer == 79)
||(x_pointer == 71 && y_pointer == 79)
||(x_pointer == 72 && y_pointer == 79)
||(x_pointer == 73 && y_pointer == 79)
||(x_pointer == 74 && y_pointer == 79)
||(x_pointer == 75 && y_pointer == 79)
||(x_pointer == 76 && y_pointer == 79)
||(x_pointer == 77 && y_pointer == 79)
||(x_pointer == 78 && y_pointer == 79)
||(x_pointer == 79 && y_pointer == 79)
||(x_pointer == 80 && y_pointer == 79)
||(x_pointer == 81 && y_pointer == 79)
||(x_pointer == 82 && y_pointer == 79)
||(x_pointer == 83 && y_pointer == 79)
||(x_pointer == 84 && y_pointer == 79)
||(x_pointer == 85 && y_pointer == 79)
||(x_pointer == 86 && y_pointer == 79)
||(x_pointer == 87 && y_pointer == 79)
||(x_pointer == 88 && y_pointer == 79)
||(x_pointer == 89 && y_pointer == 79)
||(x_pointer == 90 && y_pointer == 79)
||(x_pointer == 91 && y_pointer == 79)
||(x_pointer == 92 && y_pointer == 79)
||(x_pointer == 93 && y_pointer == 79)
||(x_pointer == 94 && y_pointer == 79)
||(x_pointer == 95 && y_pointer == 79)
||(x_pointer == 96 && y_pointer == 79)
||(x_pointer == 97 && y_pointer == 79)
||(x_pointer == 98 && y_pointer == 79)
||(x_pointer == 99 && y_pointer == 79)
||(x_pointer == 100 && y_pointer == 79)
||(x_pointer == 101 && y_pointer == 79)
||(x_pointer == 102 && y_pointer == 79)
||(x_pointer == 103 && y_pointer == 79)
||(x_pointer == 104 && y_pointer == 79)
||(x_pointer == 105 && y_pointer == 79)
||(x_pointer == 106 && y_pointer == 79)
||(x_pointer == 155 && y_pointer == 79)
||(x_pointer == 156 && y_pointer == 79)
||(x_pointer == 157 && y_pointer == 79)
||(x_pointer == 2 && y_pointer == 80)
||(x_pointer == 3 && y_pointer == 80)
||(x_pointer == 4 && y_pointer == 80)
||(x_pointer == 56 && y_pointer == 80)
||(x_pointer == 57 && y_pointer == 80)
||(x_pointer == 58 && y_pointer == 80)
||(x_pointer == 59 && y_pointer == 80)
||(x_pointer == 60 && y_pointer == 80)
||(x_pointer == 61 && y_pointer == 80)
||(x_pointer == 62 && y_pointer == 80)
||(x_pointer == 63 && y_pointer == 80)
||(x_pointer == 64 && y_pointer == 80)
||(x_pointer == 65 && y_pointer == 80)
||(x_pointer == 66 && y_pointer == 80)
||(x_pointer == 67 && y_pointer == 80)
||(x_pointer == 68 && y_pointer == 80)
||(x_pointer == 69 && y_pointer == 80)
||(x_pointer == 70 && y_pointer == 80)
||(x_pointer == 71 && y_pointer == 80)
||(x_pointer == 72 && y_pointer == 80)
||(x_pointer == 73 && y_pointer == 80)
||(x_pointer == 74 && y_pointer == 80)
||(x_pointer == 75 && y_pointer == 80)
||(x_pointer == 76 && y_pointer == 80)
||(x_pointer == 77 && y_pointer == 80)
||(x_pointer == 78 && y_pointer == 80)
||(x_pointer == 79 && y_pointer == 80)
||(x_pointer == 80 && y_pointer == 80)
||(x_pointer == 81 && y_pointer == 80)
||(x_pointer == 82 && y_pointer == 80)
||(x_pointer == 83 && y_pointer == 80)
||(x_pointer == 84 && y_pointer == 80)
||(x_pointer == 85 && y_pointer == 80)
||(x_pointer == 86 && y_pointer == 80)
||(x_pointer == 87 && y_pointer == 80)
||(x_pointer == 88 && y_pointer == 80)
||(x_pointer == 89 && y_pointer == 80)
||(x_pointer == 90 && y_pointer == 80)
||(x_pointer == 91 && y_pointer == 80)
||(x_pointer == 92 && y_pointer == 80)
||(x_pointer == 93 && y_pointer == 80)
||(x_pointer == 94 && y_pointer == 80)
||(x_pointer == 95 && y_pointer == 80)
||(x_pointer == 96 && y_pointer == 80)
||(x_pointer == 97 && y_pointer == 80)
||(x_pointer == 98 && y_pointer == 80)
||(x_pointer == 99 && y_pointer == 80)
||(x_pointer == 100 && y_pointer == 80)
||(x_pointer == 101 && y_pointer == 80)
||(x_pointer == 102 && y_pointer == 80)
||(x_pointer == 103 && y_pointer == 80)
||(x_pointer == 104 && y_pointer == 80)
||(x_pointer == 105 && y_pointer == 80)
||(x_pointer == 106 && y_pointer == 80)
||(x_pointer == 155 && y_pointer == 80)
||(x_pointer == 156 && y_pointer == 80)
||(x_pointer == 157 && y_pointer == 80)
||(x_pointer == 2 && y_pointer == 81)
||(x_pointer == 3 && y_pointer == 81)
||(x_pointer == 4 && y_pointer == 81)
||(x_pointer == 56 && y_pointer == 81)
||(x_pointer == 57 && y_pointer == 81)
||(x_pointer == 58 && y_pointer == 81)
||(x_pointer == 59 && y_pointer == 81)
||(x_pointer == 60 && y_pointer == 81)
||(x_pointer == 61 && y_pointer == 81)
||(x_pointer == 62 && y_pointer == 81)
||(x_pointer == 63 && y_pointer == 81)
||(x_pointer == 64 && y_pointer == 81)
||(x_pointer == 65 && y_pointer == 81)
||(x_pointer == 66 && y_pointer == 81)
||(x_pointer == 67 && y_pointer == 81)
||(x_pointer == 68 && y_pointer == 81)
||(x_pointer == 69 && y_pointer == 81)
||(x_pointer == 70 && y_pointer == 81)
||(x_pointer == 71 && y_pointer == 81)
||(x_pointer == 72 && y_pointer == 81)
||(x_pointer == 73 && y_pointer == 81)
||(x_pointer == 74 && y_pointer == 81)
||(x_pointer == 75 && y_pointer == 81)
||(x_pointer == 76 && y_pointer == 81)
||(x_pointer == 77 && y_pointer == 81)
||(x_pointer == 78 && y_pointer == 81)
||(x_pointer == 79 && y_pointer == 81)
||(x_pointer == 80 && y_pointer == 81)
||(x_pointer == 81 && y_pointer == 81)
||(x_pointer == 82 && y_pointer == 81)
||(x_pointer == 83 && y_pointer == 81)
||(x_pointer == 84 && y_pointer == 81)
||(x_pointer == 85 && y_pointer == 81)
||(x_pointer == 86 && y_pointer == 81)
||(x_pointer == 87 && y_pointer == 81)
||(x_pointer == 88 && y_pointer == 81)
||(x_pointer == 89 && y_pointer == 81)
||(x_pointer == 90 && y_pointer == 81)
||(x_pointer == 91 && y_pointer == 81)
||(x_pointer == 92 && y_pointer == 81)
||(x_pointer == 93 && y_pointer == 81)
||(x_pointer == 94 && y_pointer == 81)
||(x_pointer == 95 && y_pointer == 81)
||(x_pointer == 96 && y_pointer == 81)
||(x_pointer == 97 && y_pointer == 81)
||(x_pointer == 98 && y_pointer == 81)
||(x_pointer == 99 && y_pointer == 81)
||(x_pointer == 100 && y_pointer == 81)
||(x_pointer == 101 && y_pointer == 81)
||(x_pointer == 102 && y_pointer == 81)
||(x_pointer == 103 && y_pointer == 81)
||(x_pointer == 104 && y_pointer == 81)
||(x_pointer == 105 && y_pointer == 81)
||(x_pointer == 106 && y_pointer == 81)
||(x_pointer == 155 && y_pointer == 81)
||(x_pointer == 156 && y_pointer == 81)
||(x_pointer == 157 && y_pointer == 81)
||(x_pointer == 2 && y_pointer == 82)
||(x_pointer == 3 && y_pointer == 82)
||(x_pointer == 4 && y_pointer == 82)
||(x_pointer == 56 && y_pointer == 82)
||(x_pointer == 57 && y_pointer == 82)
||(x_pointer == 58 && y_pointer == 82)
||(x_pointer == 59 && y_pointer == 82)
||(x_pointer == 60 && y_pointer == 82)
||(x_pointer == 61 && y_pointer == 82)
||(x_pointer == 62 && y_pointer == 82)
||(x_pointer == 63 && y_pointer == 82)
||(x_pointer == 64 && y_pointer == 82)
||(x_pointer == 65 && y_pointer == 82)
||(x_pointer == 66 && y_pointer == 82)
||(x_pointer == 67 && y_pointer == 82)
||(x_pointer == 68 && y_pointer == 82)
||(x_pointer == 69 && y_pointer == 82)
||(x_pointer == 70 && y_pointer == 82)
||(x_pointer == 71 && y_pointer == 82)
||(x_pointer == 72 && y_pointer == 82)
||(x_pointer == 73 && y_pointer == 82)
||(x_pointer == 74 && y_pointer == 82)
||(x_pointer == 75 && y_pointer == 82)
||(x_pointer == 76 && y_pointer == 82)
||(x_pointer == 77 && y_pointer == 82)
||(x_pointer == 78 && y_pointer == 82)
||(x_pointer == 79 && y_pointer == 82)
||(x_pointer == 80 && y_pointer == 82)
||(x_pointer == 81 && y_pointer == 82)
||(x_pointer == 82 && y_pointer == 82)
||(x_pointer == 83 && y_pointer == 82)
||(x_pointer == 84 && y_pointer == 82)
||(x_pointer == 85 && y_pointer == 82)
||(x_pointer == 86 && y_pointer == 82)
||(x_pointer == 87 && y_pointer == 82)
||(x_pointer == 88 && y_pointer == 82)
||(x_pointer == 89 && y_pointer == 82)
||(x_pointer == 90 && y_pointer == 82)
||(x_pointer == 91 && y_pointer == 82)
||(x_pointer == 92 && y_pointer == 82)
||(x_pointer == 93 && y_pointer == 82)
||(x_pointer == 94 && y_pointer == 82)
||(x_pointer == 95 && y_pointer == 82)
||(x_pointer == 96 && y_pointer == 82)
||(x_pointer == 97 && y_pointer == 82)
||(x_pointer == 98 && y_pointer == 82)
||(x_pointer == 99 && y_pointer == 82)
||(x_pointer == 100 && y_pointer == 82)
||(x_pointer == 101 && y_pointer == 82)
||(x_pointer == 102 && y_pointer == 82)
||(x_pointer == 103 && y_pointer == 82)
||(x_pointer == 104 && y_pointer == 82)
||(x_pointer == 105 && y_pointer == 82)
||(x_pointer == 106 && y_pointer == 82)
||(x_pointer == 155 && y_pointer == 82)
||(x_pointer == 156 && y_pointer == 82)
||(x_pointer == 157 && y_pointer == 82)
||(x_pointer == 2 && y_pointer == 83)
||(x_pointer == 3 && y_pointer == 83)
||(x_pointer == 4 && y_pointer == 83)
||(x_pointer == 56 && y_pointer == 83)
||(x_pointer == 57 && y_pointer == 83)
||(x_pointer == 58 && y_pointer == 83)
||(x_pointer == 59 && y_pointer == 83)
||(x_pointer == 60 && y_pointer == 83)
||(x_pointer == 61 && y_pointer == 83)
||(x_pointer == 62 && y_pointer == 83)
||(x_pointer == 63 && y_pointer == 83)
||(x_pointer == 64 && y_pointer == 83)
||(x_pointer == 65 && y_pointer == 83)
||(x_pointer == 66 && y_pointer == 83)
||(x_pointer == 67 && y_pointer == 83)
||(x_pointer == 68 && y_pointer == 83)
||(x_pointer == 69 && y_pointer == 83)
||(x_pointer == 70 && y_pointer == 83)
||(x_pointer == 71 && y_pointer == 83)
||(x_pointer == 72 && y_pointer == 83)
||(x_pointer == 73 && y_pointer == 83)
||(x_pointer == 74 && y_pointer == 83)
||(x_pointer == 75 && y_pointer == 83)
||(x_pointer == 76 && y_pointer == 83)
||(x_pointer == 77 && y_pointer == 83)
||(x_pointer == 78 && y_pointer == 83)
||(x_pointer == 79 && y_pointer == 83)
||(x_pointer == 80 && y_pointer == 83)
||(x_pointer == 81 && y_pointer == 83)
||(x_pointer == 82 && y_pointer == 83)
||(x_pointer == 83 && y_pointer == 83)
||(x_pointer == 84 && y_pointer == 83)
||(x_pointer == 85 && y_pointer == 83)
||(x_pointer == 86 && y_pointer == 83)
||(x_pointer == 87 && y_pointer == 83)
||(x_pointer == 88 && y_pointer == 83)
||(x_pointer == 89 && y_pointer == 83)
||(x_pointer == 90 && y_pointer == 83)
||(x_pointer == 91 && y_pointer == 83)
||(x_pointer == 92 && y_pointer == 83)
||(x_pointer == 93 && y_pointer == 83)
||(x_pointer == 94 && y_pointer == 83)
||(x_pointer == 95 && y_pointer == 83)
||(x_pointer == 96 && y_pointer == 83)
||(x_pointer == 97 && y_pointer == 83)
||(x_pointer == 98 && y_pointer == 83)
||(x_pointer == 99 && y_pointer == 83)
||(x_pointer == 100 && y_pointer == 83)
||(x_pointer == 101 && y_pointer == 83)
||(x_pointer == 102 && y_pointer == 83)
||(x_pointer == 103 && y_pointer == 83)
||(x_pointer == 104 && y_pointer == 83)
||(x_pointer == 105 && y_pointer == 83)
||(x_pointer == 106 && y_pointer == 83)
||(x_pointer == 155 && y_pointer == 83)
||(x_pointer == 156 && y_pointer == 83)
||(x_pointer == 157 && y_pointer == 83)
||(x_pointer == 2 && y_pointer == 84)
||(x_pointer == 3 && y_pointer == 84)
||(x_pointer == 4 && y_pointer == 84)
||(x_pointer == 56 && y_pointer == 84)
||(x_pointer == 57 && y_pointer == 84)
||(x_pointer == 58 && y_pointer == 84)
||(x_pointer == 59 && y_pointer == 84)
||(x_pointer == 60 && y_pointer == 84)
||(x_pointer == 61 && y_pointer == 84)
||(x_pointer == 62 && y_pointer == 84)
||(x_pointer == 63 && y_pointer == 84)
||(x_pointer == 64 && y_pointer == 84)
||(x_pointer == 65 && y_pointer == 84)
||(x_pointer == 66 && y_pointer == 84)
||(x_pointer == 67 && y_pointer == 84)
||(x_pointer == 68 && y_pointer == 84)
||(x_pointer == 69 && y_pointer == 84)
||(x_pointer == 70 && y_pointer == 84)
||(x_pointer == 92 && y_pointer == 84)
||(x_pointer == 93 && y_pointer == 84)
||(x_pointer == 94 && y_pointer == 84)
||(x_pointer == 95 && y_pointer == 84)
||(x_pointer == 96 && y_pointer == 84)
||(x_pointer == 97 && y_pointer == 84)
||(x_pointer == 98 && y_pointer == 84)
||(x_pointer == 99 && y_pointer == 84)
||(x_pointer == 100 && y_pointer == 84)
||(x_pointer == 101 && y_pointer == 84)
||(x_pointer == 102 && y_pointer == 84)
||(x_pointer == 103 && y_pointer == 84)
||(x_pointer == 104 && y_pointer == 84)
||(x_pointer == 105 && y_pointer == 84)
||(x_pointer == 106 && y_pointer == 84)
||(x_pointer == 155 && y_pointer == 84)
||(x_pointer == 156 && y_pointer == 84)
||(x_pointer == 157 && y_pointer == 84)
||(x_pointer == 2 && y_pointer == 85)
||(x_pointer == 3 && y_pointer == 85)
||(x_pointer == 4 && y_pointer == 85)
||(x_pointer == 56 && y_pointer == 85)
||(x_pointer == 57 && y_pointer == 85)
||(x_pointer == 58 && y_pointer == 85)
||(x_pointer == 59 && y_pointer == 85)
||(x_pointer == 60 && y_pointer == 85)
||(x_pointer == 61 && y_pointer == 85)
||(x_pointer == 62 && y_pointer == 85)
||(x_pointer == 63 && y_pointer == 85)
||(x_pointer == 64 && y_pointer == 85)
||(x_pointer == 65 && y_pointer == 85)
||(x_pointer == 66 && y_pointer == 85)
||(x_pointer == 67 && y_pointer == 85)
||(x_pointer == 68 && y_pointer == 85)
||(x_pointer == 69 && y_pointer == 85)
||(x_pointer == 70 && y_pointer == 85)
||(x_pointer == 92 && y_pointer == 85)
||(x_pointer == 93 && y_pointer == 85)
||(x_pointer == 94 && y_pointer == 85)
||(x_pointer == 95 && y_pointer == 85)
||(x_pointer == 96 && y_pointer == 85)
||(x_pointer == 97 && y_pointer == 85)
||(x_pointer == 98 && y_pointer == 85)
||(x_pointer == 99 && y_pointer == 85)
||(x_pointer == 100 && y_pointer == 85)
||(x_pointer == 101 && y_pointer == 85)
||(x_pointer == 102 && y_pointer == 85)
||(x_pointer == 103 && y_pointer == 85)
||(x_pointer == 104 && y_pointer == 85)
||(x_pointer == 105 && y_pointer == 85)
||(x_pointer == 106 && y_pointer == 85)
||(x_pointer == 155 && y_pointer == 85)
||(x_pointer == 156 && y_pointer == 85)
||(x_pointer == 157 && y_pointer == 85)
||(x_pointer == 2 && y_pointer == 86)
||(x_pointer == 3 && y_pointer == 86)
||(x_pointer == 4 && y_pointer == 86)
||(x_pointer == 56 && y_pointer == 86)
||(x_pointer == 57 && y_pointer == 86)
||(x_pointer == 58 && y_pointer == 86)
||(x_pointer == 59 && y_pointer == 86)
||(x_pointer == 60 && y_pointer == 86)
||(x_pointer == 61 && y_pointer == 86)
||(x_pointer == 62 && y_pointer == 86)
||(x_pointer == 63 && y_pointer == 86)
||(x_pointer == 64 && y_pointer == 86)
||(x_pointer == 65 && y_pointer == 86)
||(x_pointer == 66 && y_pointer == 86)
||(x_pointer == 67 && y_pointer == 86)
||(x_pointer == 68 && y_pointer == 86)
||(x_pointer == 69 && y_pointer == 86)
||(x_pointer == 70 && y_pointer == 86)
||(x_pointer == 92 && y_pointer == 86)
||(x_pointer == 93 && y_pointer == 86)
||(x_pointer == 94 && y_pointer == 86)
||(x_pointer == 95 && y_pointer == 86)
||(x_pointer == 96 && y_pointer == 86)
||(x_pointer == 97 && y_pointer == 86)
||(x_pointer == 98 && y_pointer == 86)
||(x_pointer == 99 && y_pointer == 86)
||(x_pointer == 100 && y_pointer == 86)
||(x_pointer == 101 && y_pointer == 86)
||(x_pointer == 102 && y_pointer == 86)
||(x_pointer == 103 && y_pointer == 86)
||(x_pointer == 104 && y_pointer == 86)
||(x_pointer == 105 && y_pointer == 86)
||(x_pointer == 106 && y_pointer == 86)
||(x_pointer == 155 && y_pointer == 86)
||(x_pointer == 156 && y_pointer == 86)
||(x_pointer == 157 && y_pointer == 86)
||(x_pointer == 2 && y_pointer == 87)
||(x_pointer == 3 && y_pointer == 87)
||(x_pointer == 4 && y_pointer == 87)
||(x_pointer == 56 && y_pointer == 87)
||(x_pointer == 57 && y_pointer == 87)
||(x_pointer == 58 && y_pointer == 87)
||(x_pointer == 59 && y_pointer == 87)
||(x_pointer == 60 && y_pointer == 87)
||(x_pointer == 61 && y_pointer == 87)
||(x_pointer == 62 && y_pointer == 87)
||(x_pointer == 63 && y_pointer == 87)
||(x_pointer == 64 && y_pointer == 87)
||(x_pointer == 65 && y_pointer == 87)
||(x_pointer == 66 && y_pointer == 87)
||(x_pointer == 67 && y_pointer == 87)
||(x_pointer == 68 && y_pointer == 87)
||(x_pointer == 69 && y_pointer == 87)
||(x_pointer == 70 && y_pointer == 87)
||(x_pointer == 92 && y_pointer == 87)
||(x_pointer == 93 && y_pointer == 87)
||(x_pointer == 94 && y_pointer == 87)
||(x_pointer == 95 && y_pointer == 87)
||(x_pointer == 96 && y_pointer == 87)
||(x_pointer == 97 && y_pointer == 87)
||(x_pointer == 98 && y_pointer == 87)
||(x_pointer == 99 && y_pointer == 87)
||(x_pointer == 100 && y_pointer == 87)
||(x_pointer == 101 && y_pointer == 87)
||(x_pointer == 102 && y_pointer == 87)
||(x_pointer == 103 && y_pointer == 87)
||(x_pointer == 104 && y_pointer == 87)
||(x_pointer == 105 && y_pointer == 87)
||(x_pointer == 106 && y_pointer == 87)
||(x_pointer == 155 && y_pointer == 87)
||(x_pointer == 156 && y_pointer == 87)
||(x_pointer == 157 && y_pointer == 87)
||(x_pointer == 2 && y_pointer == 88)
||(x_pointer == 3 && y_pointer == 88)
||(x_pointer == 4 && y_pointer == 88)
||(x_pointer == 56 && y_pointer == 88)
||(x_pointer == 57 && y_pointer == 88)
||(x_pointer == 58 && y_pointer == 88)
||(x_pointer == 59 && y_pointer == 88)
||(x_pointer == 60 && y_pointer == 88)
||(x_pointer == 61 && y_pointer == 88)
||(x_pointer == 62 && y_pointer == 88)
||(x_pointer == 63 && y_pointer == 88)
||(x_pointer == 64 && y_pointer == 88)
||(x_pointer == 65 && y_pointer == 88)
||(x_pointer == 66 && y_pointer == 88)
||(x_pointer == 67 && y_pointer == 88)
||(x_pointer == 68 && y_pointer == 88)
||(x_pointer == 69 && y_pointer == 88)
||(x_pointer == 70 && y_pointer == 88)
||(x_pointer == 92 && y_pointer == 88)
||(x_pointer == 93 && y_pointer == 88)
||(x_pointer == 94 && y_pointer == 88)
||(x_pointer == 95 && y_pointer == 88)
||(x_pointer == 96 && y_pointer == 88)
||(x_pointer == 97 && y_pointer == 88)
||(x_pointer == 98 && y_pointer == 88)
||(x_pointer == 99 && y_pointer == 88)
||(x_pointer == 100 && y_pointer == 88)
||(x_pointer == 101 && y_pointer == 88)
||(x_pointer == 102 && y_pointer == 88)
||(x_pointer == 103 && y_pointer == 88)
||(x_pointer == 104 && y_pointer == 88)
||(x_pointer == 105 && y_pointer == 88)
||(x_pointer == 106 && y_pointer == 88)
||(x_pointer == 155 && y_pointer == 88)
||(x_pointer == 156 && y_pointer == 88)
||(x_pointer == 157 && y_pointer == 88)
||(x_pointer == 2 && y_pointer == 89)
||(x_pointer == 3 && y_pointer == 89)
||(x_pointer == 4 && y_pointer == 89)
||(x_pointer == 56 && y_pointer == 89)
||(x_pointer == 57 && y_pointer == 89)
||(x_pointer == 58 && y_pointer == 89)
||(x_pointer == 59 && y_pointer == 89)
||(x_pointer == 60 && y_pointer == 89)
||(x_pointer == 61 && y_pointer == 89)
||(x_pointer == 62 && y_pointer == 89)
||(x_pointer == 63 && y_pointer == 89)
||(x_pointer == 64 && y_pointer == 89)
||(x_pointer == 65 && y_pointer == 89)
||(x_pointer == 66 && y_pointer == 89)
||(x_pointer == 67 && y_pointer == 89)
||(x_pointer == 68 && y_pointer == 89)
||(x_pointer == 69 && y_pointer == 89)
||(x_pointer == 70 && y_pointer == 89)
||(x_pointer == 92 && y_pointer == 89)
||(x_pointer == 93 && y_pointer == 89)
||(x_pointer == 94 && y_pointer == 89)
||(x_pointer == 95 && y_pointer == 89)
||(x_pointer == 96 && y_pointer == 89)
||(x_pointer == 97 && y_pointer == 89)
||(x_pointer == 98 && y_pointer == 89)
||(x_pointer == 99 && y_pointer == 89)
||(x_pointer == 100 && y_pointer == 89)
||(x_pointer == 101 && y_pointer == 89)
||(x_pointer == 102 && y_pointer == 89)
||(x_pointer == 103 && y_pointer == 89)
||(x_pointer == 104 && y_pointer == 89)
||(x_pointer == 105 && y_pointer == 89)
||(x_pointer == 106 && y_pointer == 89)
||(x_pointer == 155 && y_pointer == 89)
||(x_pointer == 156 && y_pointer == 89)
||(x_pointer == 157 && y_pointer == 89)
||(x_pointer == 2 && y_pointer == 90)
||(x_pointer == 3 && y_pointer == 90)
||(x_pointer == 4 && y_pointer == 90)
||(x_pointer == 56 && y_pointer == 90)
||(x_pointer == 57 && y_pointer == 90)
||(x_pointer == 58 && y_pointer == 90)
||(x_pointer == 59 && y_pointer == 90)
||(x_pointer == 60 && y_pointer == 90)
||(x_pointer == 61 && y_pointer == 90)
||(x_pointer == 62 && y_pointer == 90)
||(x_pointer == 63 && y_pointer == 90)
||(x_pointer == 64 && y_pointer == 90)
||(x_pointer == 65 && y_pointer == 90)
||(x_pointer == 66 && y_pointer == 90)
||(x_pointer == 67 && y_pointer == 90)
||(x_pointer == 68 && y_pointer == 90)
||(x_pointer == 69 && y_pointer == 90)
||(x_pointer == 70 && y_pointer == 90)
||(x_pointer == 92 && y_pointer == 90)
||(x_pointer == 93 && y_pointer == 90)
||(x_pointer == 94 && y_pointer == 90)
||(x_pointer == 95 && y_pointer == 90)
||(x_pointer == 96 && y_pointer == 90)
||(x_pointer == 97 && y_pointer == 90)
||(x_pointer == 98 && y_pointer == 90)
||(x_pointer == 99 && y_pointer == 90)
||(x_pointer == 100 && y_pointer == 90)
||(x_pointer == 101 && y_pointer == 90)
||(x_pointer == 102 && y_pointer == 90)
||(x_pointer == 103 && y_pointer == 90)
||(x_pointer == 104 && y_pointer == 90)
||(x_pointer == 105 && y_pointer == 90)
||(x_pointer == 106 && y_pointer == 90)
||(x_pointer == 155 && y_pointer == 90)
||(x_pointer == 156 && y_pointer == 90)
||(x_pointer == 157 && y_pointer == 90)
||(x_pointer == 2 && y_pointer == 91)
||(x_pointer == 3 && y_pointer == 91)
||(x_pointer == 4 && y_pointer == 91)
||(x_pointer == 56 && y_pointer == 91)
||(x_pointer == 57 && y_pointer == 91)
||(x_pointer == 58 && y_pointer == 91)
||(x_pointer == 59 && y_pointer == 91)
||(x_pointer == 60 && y_pointer == 91)
||(x_pointer == 61 && y_pointer == 91)
||(x_pointer == 62 && y_pointer == 91)
||(x_pointer == 63 && y_pointer == 91)
||(x_pointer == 64 && y_pointer == 91)
||(x_pointer == 65 && y_pointer == 91)
||(x_pointer == 66 && y_pointer == 91)
||(x_pointer == 67 && y_pointer == 91)
||(x_pointer == 68 && y_pointer == 91)
||(x_pointer == 69 && y_pointer == 91)
||(x_pointer == 70 && y_pointer == 91)
||(x_pointer == 92 && y_pointer == 91)
||(x_pointer == 93 && y_pointer == 91)
||(x_pointer == 94 && y_pointer == 91)
||(x_pointer == 95 && y_pointer == 91)
||(x_pointer == 96 && y_pointer == 91)
||(x_pointer == 97 && y_pointer == 91)
||(x_pointer == 98 && y_pointer == 91)
||(x_pointer == 99 && y_pointer == 91)
||(x_pointer == 100 && y_pointer == 91)
||(x_pointer == 101 && y_pointer == 91)
||(x_pointer == 102 && y_pointer == 91)
||(x_pointer == 103 && y_pointer == 91)
||(x_pointer == 104 && y_pointer == 91)
||(x_pointer == 105 && y_pointer == 91)
||(x_pointer == 106 && y_pointer == 91)
||(x_pointer == 155 && y_pointer == 91)
||(x_pointer == 156 && y_pointer == 91)
||(x_pointer == 157 && y_pointer == 91)
||(x_pointer == 2 && y_pointer == 92)
||(x_pointer == 3 && y_pointer == 92)
||(x_pointer == 4 && y_pointer == 92)
||(x_pointer == 56 && y_pointer == 92)
||(x_pointer == 57 && y_pointer == 92)
||(x_pointer == 58 && y_pointer == 92)
||(x_pointer == 59 && y_pointer == 92)
||(x_pointer == 60 && y_pointer == 92)
||(x_pointer == 61 && y_pointer == 92)
||(x_pointer == 62 && y_pointer == 92)
||(x_pointer == 63 && y_pointer == 92)
||(x_pointer == 64 && y_pointer == 92)
||(x_pointer == 65 && y_pointer == 92)
||(x_pointer == 66 && y_pointer == 92)
||(x_pointer == 67 && y_pointer == 92)
||(x_pointer == 68 && y_pointer == 92)
||(x_pointer == 69 && y_pointer == 92)
||(x_pointer == 70 && y_pointer == 92)
||(x_pointer == 92 && y_pointer == 92)
||(x_pointer == 93 && y_pointer == 92)
||(x_pointer == 94 && y_pointer == 92)
||(x_pointer == 95 && y_pointer == 92)
||(x_pointer == 96 && y_pointer == 92)
||(x_pointer == 97 && y_pointer == 92)
||(x_pointer == 98 && y_pointer == 92)
||(x_pointer == 99 && y_pointer == 92)
||(x_pointer == 100 && y_pointer == 92)
||(x_pointer == 101 && y_pointer == 92)
||(x_pointer == 102 && y_pointer == 92)
||(x_pointer == 103 && y_pointer == 92)
||(x_pointer == 104 && y_pointer == 92)
||(x_pointer == 105 && y_pointer == 92)
||(x_pointer == 106 && y_pointer == 92)
||(x_pointer == 155 && y_pointer == 92)
||(x_pointer == 156 && y_pointer == 92)
||(x_pointer == 157 && y_pointer == 92)
||(x_pointer == 2 && y_pointer == 93)
||(x_pointer == 3 && y_pointer == 93)
||(x_pointer == 4 && y_pointer == 93)
||(x_pointer == 56 && y_pointer == 93)
||(x_pointer == 57 && y_pointer == 93)
||(x_pointer == 58 && y_pointer == 93)
||(x_pointer == 59 && y_pointer == 93)
||(x_pointer == 60 && y_pointer == 93)
||(x_pointer == 61 && y_pointer == 93)
||(x_pointer == 62 && y_pointer == 93)
||(x_pointer == 63 && y_pointer == 93)
||(x_pointer == 64 && y_pointer == 93)
||(x_pointer == 65 && y_pointer == 93)
||(x_pointer == 66 && y_pointer == 93)
||(x_pointer == 67 && y_pointer == 93)
||(x_pointer == 68 && y_pointer == 93)
||(x_pointer == 69 && y_pointer == 93)
||(x_pointer == 70 && y_pointer == 93)
||(x_pointer == 92 && y_pointer == 93)
||(x_pointer == 93 && y_pointer == 93)
||(x_pointer == 94 && y_pointer == 93)
||(x_pointer == 95 && y_pointer == 93)
||(x_pointer == 96 && y_pointer == 93)
||(x_pointer == 97 && y_pointer == 93)
||(x_pointer == 98 && y_pointer == 93)
||(x_pointer == 99 && y_pointer == 93)
||(x_pointer == 100 && y_pointer == 93)
||(x_pointer == 101 && y_pointer == 93)
||(x_pointer == 102 && y_pointer == 93)
||(x_pointer == 103 && y_pointer == 93)
||(x_pointer == 104 && y_pointer == 93)
||(x_pointer == 105 && y_pointer == 93)
||(x_pointer == 106 && y_pointer == 93)
||(x_pointer == 155 && y_pointer == 93)
||(x_pointer == 156 && y_pointer == 93)
||(x_pointer == 157 && y_pointer == 93)
||(x_pointer == 2 && y_pointer == 94)
||(x_pointer == 3 && y_pointer == 94)
||(x_pointer == 4 && y_pointer == 94)
||(x_pointer == 56 && y_pointer == 94)
||(x_pointer == 57 && y_pointer == 94)
||(x_pointer == 58 && y_pointer == 94)
||(x_pointer == 59 && y_pointer == 94)
||(x_pointer == 60 && y_pointer == 94)
||(x_pointer == 61 && y_pointer == 94)
||(x_pointer == 62 && y_pointer == 94)
||(x_pointer == 63 && y_pointer == 94)
||(x_pointer == 64 && y_pointer == 94)
||(x_pointer == 65 && y_pointer == 94)
||(x_pointer == 66 && y_pointer == 94)
||(x_pointer == 67 && y_pointer == 94)
||(x_pointer == 68 && y_pointer == 94)
||(x_pointer == 69 && y_pointer == 94)
||(x_pointer == 70 && y_pointer == 94)
||(x_pointer == 92 && y_pointer == 94)
||(x_pointer == 93 && y_pointer == 94)
||(x_pointer == 94 && y_pointer == 94)
||(x_pointer == 95 && y_pointer == 94)
||(x_pointer == 96 && y_pointer == 94)
||(x_pointer == 97 && y_pointer == 94)
||(x_pointer == 98 && y_pointer == 94)
||(x_pointer == 99 && y_pointer == 94)
||(x_pointer == 100 && y_pointer == 94)
||(x_pointer == 101 && y_pointer == 94)
||(x_pointer == 102 && y_pointer == 94)
||(x_pointer == 103 && y_pointer == 94)
||(x_pointer == 104 && y_pointer == 94)
||(x_pointer == 105 && y_pointer == 94)
||(x_pointer == 106 && y_pointer == 94)
||(x_pointer == 155 && y_pointer == 94)
||(x_pointer == 156 && y_pointer == 94)
||(x_pointer == 157 && y_pointer == 94)
||(x_pointer == 2 && y_pointer == 95)
||(x_pointer == 3 && y_pointer == 95)
||(x_pointer == 4 && y_pointer == 95)
||(x_pointer == 56 && y_pointer == 95)
||(x_pointer == 57 && y_pointer == 95)
||(x_pointer == 58 && y_pointer == 95)
||(x_pointer == 59 && y_pointer == 95)
||(x_pointer == 60 && y_pointer == 95)
||(x_pointer == 61 && y_pointer == 95)
||(x_pointer == 62 && y_pointer == 95)
||(x_pointer == 63 && y_pointer == 95)
||(x_pointer == 64 && y_pointer == 95)
||(x_pointer == 65 && y_pointer == 95)
||(x_pointer == 66 && y_pointer == 95)
||(x_pointer == 67 && y_pointer == 95)
||(x_pointer == 68 && y_pointer == 95)
||(x_pointer == 69 && y_pointer == 95)
||(x_pointer == 70 && y_pointer == 95)
||(x_pointer == 92 && y_pointer == 95)
||(x_pointer == 93 && y_pointer == 95)
||(x_pointer == 94 && y_pointer == 95)
||(x_pointer == 95 && y_pointer == 95)
||(x_pointer == 96 && y_pointer == 95)
||(x_pointer == 97 && y_pointer == 95)
||(x_pointer == 98 && y_pointer == 95)
||(x_pointer == 99 && y_pointer == 95)
||(x_pointer == 100 && y_pointer == 95)
||(x_pointer == 101 && y_pointer == 95)
||(x_pointer == 102 && y_pointer == 95)
||(x_pointer == 103 && y_pointer == 95)
||(x_pointer == 104 && y_pointer == 95)
||(x_pointer == 105 && y_pointer == 95)
||(x_pointer == 106 && y_pointer == 95)
||(x_pointer == 155 && y_pointer == 95)
||(x_pointer == 156 && y_pointer == 95)
||(x_pointer == 157 && y_pointer == 95)
||(x_pointer == 2 && y_pointer == 96)
||(x_pointer == 3 && y_pointer == 96)
||(x_pointer == 4 && y_pointer == 96)
||(x_pointer == 56 && y_pointer == 96)
||(x_pointer == 57 && y_pointer == 96)
||(x_pointer == 58 && y_pointer == 96)
||(x_pointer == 59 && y_pointer == 96)
||(x_pointer == 60 && y_pointer == 96)
||(x_pointer == 61 && y_pointer == 96)
||(x_pointer == 62 && y_pointer == 96)
||(x_pointer == 63 && y_pointer == 96)
||(x_pointer == 64 && y_pointer == 96)
||(x_pointer == 65 && y_pointer == 96)
||(x_pointer == 66 && y_pointer == 96)
||(x_pointer == 67 && y_pointer == 96)
||(x_pointer == 68 && y_pointer == 96)
||(x_pointer == 69 && y_pointer == 96)
||(x_pointer == 70 && y_pointer == 96)
||(x_pointer == 92 && y_pointer == 96)
||(x_pointer == 93 && y_pointer == 96)
||(x_pointer == 94 && y_pointer == 96)
||(x_pointer == 95 && y_pointer == 96)
||(x_pointer == 96 && y_pointer == 96)
||(x_pointer == 97 && y_pointer == 96)
||(x_pointer == 98 && y_pointer == 96)
||(x_pointer == 99 && y_pointer == 96)
||(x_pointer == 100 && y_pointer == 96)
||(x_pointer == 101 && y_pointer == 96)
||(x_pointer == 102 && y_pointer == 96)
||(x_pointer == 103 && y_pointer == 96)
||(x_pointer == 104 && y_pointer == 96)
||(x_pointer == 105 && y_pointer == 96)
||(x_pointer == 106 && y_pointer == 96)
||(x_pointer == 155 && y_pointer == 96)
||(x_pointer == 156 && y_pointer == 96)
||(x_pointer == 157 && y_pointer == 96)
||(x_pointer == 2 && y_pointer == 97)
||(x_pointer == 3 && y_pointer == 97)
||(x_pointer == 4 && y_pointer == 97)
||(x_pointer == 56 && y_pointer == 97)
||(x_pointer == 57 && y_pointer == 97)
||(x_pointer == 58 && y_pointer == 97)
||(x_pointer == 59 && y_pointer == 97)
||(x_pointer == 60 && y_pointer == 97)
||(x_pointer == 61 && y_pointer == 97)
||(x_pointer == 62 && y_pointer == 97)
||(x_pointer == 63 && y_pointer == 97)
||(x_pointer == 64 && y_pointer == 97)
||(x_pointer == 65 && y_pointer == 97)
||(x_pointer == 66 && y_pointer == 97)
||(x_pointer == 67 && y_pointer == 97)
||(x_pointer == 68 && y_pointer == 97)
||(x_pointer == 69 && y_pointer == 97)
||(x_pointer == 70 && y_pointer == 97)
||(x_pointer == 92 && y_pointer == 97)
||(x_pointer == 93 && y_pointer == 97)
||(x_pointer == 94 && y_pointer == 97)
||(x_pointer == 95 && y_pointer == 97)
||(x_pointer == 96 && y_pointer == 97)
||(x_pointer == 97 && y_pointer == 97)
||(x_pointer == 98 && y_pointer == 97)
||(x_pointer == 99 && y_pointer == 97)
||(x_pointer == 100 && y_pointer == 97)
||(x_pointer == 101 && y_pointer == 97)
||(x_pointer == 102 && y_pointer == 97)
||(x_pointer == 103 && y_pointer == 97)
||(x_pointer == 104 && y_pointer == 97)
||(x_pointer == 105 && y_pointer == 97)
||(x_pointer == 106 && y_pointer == 97)
||(x_pointer == 155 && y_pointer == 97)
||(x_pointer == 156 && y_pointer == 97)
||(x_pointer == 157 && y_pointer == 97)
||(x_pointer == 2 && y_pointer == 98)
||(x_pointer == 3 && y_pointer == 98)
||(x_pointer == 4 && y_pointer == 98)
||(x_pointer == 155 && y_pointer == 98)
||(x_pointer == 156 && y_pointer == 98)
||(x_pointer == 157 && y_pointer == 98)
||(x_pointer == 2 && y_pointer == 99)
||(x_pointer == 3 && y_pointer == 99)
||(x_pointer == 4 && y_pointer == 99)
||(x_pointer == 155 && y_pointer == 99)
||(x_pointer == 156 && y_pointer == 99)
||(x_pointer == 157 && y_pointer == 99)
||(x_pointer == 2 && y_pointer == 100)
||(x_pointer == 3 && y_pointer == 100)
||(x_pointer == 4 && y_pointer == 100)
||(x_pointer == 155 && y_pointer == 100)
||(x_pointer == 156 && y_pointer == 100)
||(x_pointer == 157 && y_pointer == 100)
||(x_pointer == 2 && y_pointer == 101)
||(x_pointer == 3 && y_pointer == 101)
||(x_pointer == 4 && y_pointer == 101)
||(x_pointer == 155 && y_pointer == 101)
||(x_pointer == 156 && y_pointer == 101)
||(x_pointer == 157 && y_pointer == 101)
||(x_pointer == 2 && y_pointer == 102)
||(x_pointer == 3 && y_pointer == 102)
||(x_pointer == 4 && y_pointer == 102)
||(x_pointer == 155 && y_pointer == 102)
||(x_pointer == 156 && y_pointer == 102)
||(x_pointer == 157 && y_pointer == 102)
||(x_pointer == 2 && y_pointer == 103)
||(x_pointer == 3 && y_pointer == 103)
||(x_pointer == 4 && y_pointer == 103)
||(x_pointer == 155 && y_pointer == 103)
||(x_pointer == 156 && y_pointer == 103)
||(x_pointer == 157 && y_pointer == 103)
||(x_pointer == 2 && y_pointer == 104)
||(x_pointer == 3 && y_pointer == 104)
||(x_pointer == 4 && y_pointer == 104)
||(x_pointer == 155 && y_pointer == 104)
||(x_pointer == 156 && y_pointer == 104)
||(x_pointer == 157 && y_pointer == 104)
||(x_pointer == 2 && y_pointer == 105)
||(x_pointer == 3 && y_pointer == 105)
||(x_pointer == 4 && y_pointer == 105)
||(x_pointer == 155 && y_pointer == 105)
||(x_pointer == 156 && y_pointer == 105)
||(x_pointer == 157 && y_pointer == 105)
||(x_pointer == 2 && y_pointer == 106)
||(x_pointer == 3 && y_pointer == 106)
||(x_pointer == 4 && y_pointer == 106)
||(x_pointer == 155 && y_pointer == 106)
||(x_pointer == 156 && y_pointer == 106)
||(x_pointer == 157 && y_pointer == 106)
||(x_pointer == 2 && y_pointer == 107)
||(x_pointer == 3 && y_pointer == 107)
||(x_pointer == 4 && y_pointer == 107)
||(x_pointer == 155 && y_pointer == 107)
||(x_pointer == 156 && y_pointer == 107)
||(x_pointer == 157 && y_pointer == 107)
||(x_pointer == 2 && y_pointer == 108)
||(x_pointer == 3 && y_pointer == 108)
||(x_pointer == 4 && y_pointer == 108)
||(x_pointer == 155 && y_pointer == 108)
||(x_pointer == 156 && y_pointer == 108)
||(x_pointer == 157 && y_pointer == 108)
||(x_pointer == 2 && y_pointer == 109)
||(x_pointer == 3 && y_pointer == 109)
||(x_pointer == 4 && y_pointer == 109)
||(x_pointer == 155 && y_pointer == 109)
||(x_pointer == 156 && y_pointer == 109)
||(x_pointer == 157 && y_pointer == 109)
||(x_pointer == 2 && y_pointer == 110)
||(x_pointer == 3 && y_pointer == 110)
||(x_pointer == 4 && y_pointer == 110)
||(x_pointer == 5 && y_pointer == 110)
||(x_pointer == 6 && y_pointer == 110)
||(x_pointer == 7 && y_pointer == 110)
||(x_pointer == 8 && y_pointer == 110)
||(x_pointer == 9 && y_pointer == 110)
||(x_pointer == 10 && y_pointer == 110)
||(x_pointer == 11 && y_pointer == 110)
||(x_pointer == 12 && y_pointer == 110)
||(x_pointer == 13 && y_pointer == 110)
||(x_pointer == 14 && y_pointer == 110)
||(x_pointer == 15 && y_pointer == 110)
||(x_pointer == 16 && y_pointer == 110)
||(x_pointer == 17 && y_pointer == 110)
||(x_pointer == 18 && y_pointer == 110)
||(x_pointer == 19 && y_pointer == 110)
||(x_pointer == 20 && y_pointer == 110)
||(x_pointer == 21 && y_pointer == 110)
||(x_pointer == 22 && y_pointer == 110)
||(x_pointer == 23 && y_pointer == 110)
||(x_pointer == 24 && y_pointer == 110)
||(x_pointer == 25 && y_pointer == 110)
||(x_pointer == 26 && y_pointer == 110)
||(x_pointer == 27 && y_pointer == 110)
||(x_pointer == 28 && y_pointer == 110)
||(x_pointer == 29 && y_pointer == 110)
||(x_pointer == 30 && y_pointer == 110)
||(x_pointer == 31 && y_pointer == 110)
||(x_pointer == 32 && y_pointer == 110)
||(x_pointer == 33 && y_pointer == 110)
||(x_pointer == 34 && y_pointer == 110)
||(x_pointer == 35 && y_pointer == 110)
||(x_pointer == 36 && y_pointer == 110)
||(x_pointer == 37 && y_pointer == 110)
||(x_pointer == 38 && y_pointer == 110)
||(x_pointer == 39 && y_pointer == 110)
||(x_pointer == 40 && y_pointer == 110)
||(x_pointer == 41 && y_pointer == 110)
||(x_pointer == 42 && y_pointer == 110)
||(x_pointer == 43 && y_pointer == 110)
||(x_pointer == 44 && y_pointer == 110)
||(x_pointer == 45 && y_pointer == 110)
||(x_pointer == 46 && y_pointer == 110)
||(x_pointer == 47 && y_pointer == 110)
||(x_pointer == 48 && y_pointer == 110)
||(x_pointer == 49 && y_pointer == 110)
||(x_pointer == 50 && y_pointer == 110)
||(x_pointer == 51 && y_pointer == 110)
||(x_pointer == 52 && y_pointer == 110)
||(x_pointer == 53 && y_pointer == 110)
||(x_pointer == 54 && y_pointer == 110)
||(x_pointer == 55 && y_pointer == 110)
||(x_pointer == 56 && y_pointer == 110)
||(x_pointer == 57 && y_pointer == 110)
||(x_pointer == 58 && y_pointer == 110)
||(x_pointer == 59 && y_pointer == 110)
||(x_pointer == 60 && y_pointer == 110)
||(x_pointer == 61 && y_pointer == 110)
||(x_pointer == 62 && y_pointer == 110)
||(x_pointer == 63 && y_pointer == 110)
||(x_pointer == 64 && y_pointer == 110)
||(x_pointer == 65 && y_pointer == 110)
||(x_pointer == 66 && y_pointer == 110)
||(x_pointer == 67 && y_pointer == 110)
||(x_pointer == 68 && y_pointer == 110)
||(x_pointer == 69 && y_pointer == 110)
||(x_pointer == 70 && y_pointer == 110)
||(x_pointer == 71 && y_pointer == 110)
||(x_pointer == 72 && y_pointer == 110)
||(x_pointer == 73 && y_pointer == 110)
||(x_pointer == 74 && y_pointer == 110)
||(x_pointer == 75 && y_pointer == 110)
||(x_pointer == 76 && y_pointer == 110)
||(x_pointer == 77 && y_pointer == 110)
||(x_pointer == 78 && y_pointer == 110)
||(x_pointer == 79 && y_pointer == 110)
||(x_pointer == 80 && y_pointer == 110)
||(x_pointer == 81 && y_pointer == 110)
||(x_pointer == 82 && y_pointer == 110)
||(x_pointer == 83 && y_pointer == 110)
||(x_pointer == 84 && y_pointer == 110)
||(x_pointer == 85 && y_pointer == 110)
||(x_pointer == 86 && y_pointer == 110)
||(x_pointer == 87 && y_pointer == 110)
||(x_pointer == 88 && y_pointer == 110)
||(x_pointer == 89 && y_pointer == 110)
||(x_pointer == 90 && y_pointer == 110)
||(x_pointer == 91 && y_pointer == 110)
||(x_pointer == 92 && y_pointer == 110)
||(x_pointer == 93 && y_pointer == 110)
||(x_pointer == 94 && y_pointer == 110)
||(x_pointer == 95 && y_pointer == 110)
||(x_pointer == 96 && y_pointer == 110)
||(x_pointer == 97 && y_pointer == 110)
||(x_pointer == 98 && y_pointer == 110)
||(x_pointer == 99 && y_pointer == 110)
||(x_pointer == 100 && y_pointer == 110)
||(x_pointer == 101 && y_pointer == 110)
||(x_pointer == 102 && y_pointer == 110)
||(x_pointer == 103 && y_pointer == 110)
||(x_pointer == 104 && y_pointer == 110)
||(x_pointer == 105 && y_pointer == 110)
||(x_pointer == 106 && y_pointer == 110)
||(x_pointer == 107 && y_pointer == 110)
||(x_pointer == 108 && y_pointer == 110)
||(x_pointer == 109 && y_pointer == 110)
||(x_pointer == 110 && y_pointer == 110)
||(x_pointer == 111 && y_pointer == 110)
||(x_pointer == 112 && y_pointer == 110)
||(x_pointer == 113 && y_pointer == 110)
||(x_pointer == 114 && y_pointer == 110)
||(x_pointer == 115 && y_pointer == 110)
||(x_pointer == 116 && y_pointer == 110)
||(x_pointer == 117 && y_pointer == 110)
||(x_pointer == 118 && y_pointer == 110)
||(x_pointer == 119 && y_pointer == 110)
||(x_pointer == 120 && y_pointer == 110)
||(x_pointer == 121 && y_pointer == 110)
||(x_pointer == 122 && y_pointer == 110)
||(x_pointer == 123 && y_pointer == 110)
||(x_pointer == 124 && y_pointer == 110)
||(x_pointer == 125 && y_pointer == 110)
||(x_pointer == 126 && y_pointer == 110)
||(x_pointer == 127 && y_pointer == 110)
||(x_pointer == 128 && y_pointer == 110)
||(x_pointer == 129 && y_pointer == 110)
||(x_pointer == 130 && y_pointer == 110)
||(x_pointer == 131 && y_pointer == 110)
||(x_pointer == 132 && y_pointer == 110)
||(x_pointer == 133 && y_pointer == 110)
||(x_pointer == 134 && y_pointer == 110)
||(x_pointer == 135 && y_pointer == 110)
||(x_pointer == 136 && y_pointer == 110)
||(x_pointer == 137 && y_pointer == 110)
||(x_pointer == 138 && y_pointer == 110)
||(x_pointer == 139 && y_pointer == 110)
||(x_pointer == 140 && y_pointer == 110)
||(x_pointer == 141 && y_pointer == 110)
||(x_pointer == 142 && y_pointer == 110)
||(x_pointer == 143 && y_pointer == 110)
||(x_pointer == 144 && y_pointer == 110)
||(x_pointer == 145 && y_pointer == 110)
||(x_pointer == 146 && y_pointer == 110)
||(x_pointer == 147 && y_pointer == 110)
||(x_pointer == 148 && y_pointer == 110)
||(x_pointer == 149 && y_pointer == 110)
||(x_pointer == 150 && y_pointer == 110)
||(x_pointer == 151 && y_pointer == 110)
||(x_pointer == 152 && y_pointer == 110)
||(x_pointer == 153 && y_pointer == 110)
||(x_pointer == 154 && y_pointer == 110)
||(x_pointer == 155 && y_pointer == 110)
||(x_pointer == 156 && y_pointer == 110)
||(x_pointer == 157 && y_pointer == 110)
||(x_pointer == 2 && y_pointer == 111)
||(x_pointer == 3 && y_pointer == 111)
||(x_pointer == 4 && y_pointer == 111)
||(x_pointer == 5 && y_pointer == 111)
||(x_pointer == 6 && y_pointer == 111)
||(x_pointer == 7 && y_pointer == 111)
||(x_pointer == 8 && y_pointer == 111)
||(x_pointer == 9 && y_pointer == 111)
||(x_pointer == 10 && y_pointer == 111)
||(x_pointer == 11 && y_pointer == 111)
||(x_pointer == 12 && y_pointer == 111)
||(x_pointer == 13 && y_pointer == 111)
||(x_pointer == 14 && y_pointer == 111)
||(x_pointer == 15 && y_pointer == 111)
||(x_pointer == 16 && y_pointer == 111)
||(x_pointer == 17 && y_pointer == 111)
||(x_pointer == 18 && y_pointer == 111)
||(x_pointer == 19 && y_pointer == 111)
||(x_pointer == 20 && y_pointer == 111)
||(x_pointer == 21 && y_pointer == 111)
||(x_pointer == 22 && y_pointer == 111)
||(x_pointer == 23 && y_pointer == 111)
||(x_pointer == 24 && y_pointer == 111)
||(x_pointer == 25 && y_pointer == 111)
||(x_pointer == 26 && y_pointer == 111)
||(x_pointer == 27 && y_pointer == 111)
||(x_pointer == 28 && y_pointer == 111)
||(x_pointer == 29 && y_pointer == 111)
||(x_pointer == 30 && y_pointer == 111)
||(x_pointer == 31 && y_pointer == 111)
||(x_pointer == 32 && y_pointer == 111)
||(x_pointer == 33 && y_pointer == 111)
||(x_pointer == 34 && y_pointer == 111)
||(x_pointer == 35 && y_pointer == 111)
||(x_pointer == 36 && y_pointer == 111)
||(x_pointer == 37 && y_pointer == 111)
||(x_pointer == 38 && y_pointer == 111)
||(x_pointer == 39 && y_pointer == 111)
||(x_pointer == 40 && y_pointer == 111)
||(x_pointer == 41 && y_pointer == 111)
||(x_pointer == 42 && y_pointer == 111)
||(x_pointer == 43 && y_pointer == 111)
||(x_pointer == 44 && y_pointer == 111)
||(x_pointer == 45 && y_pointer == 111)
||(x_pointer == 46 && y_pointer == 111)
||(x_pointer == 47 && y_pointer == 111)
||(x_pointer == 48 && y_pointer == 111)
||(x_pointer == 49 && y_pointer == 111)
||(x_pointer == 50 && y_pointer == 111)
||(x_pointer == 51 && y_pointer == 111)
||(x_pointer == 52 && y_pointer == 111)
||(x_pointer == 53 && y_pointer == 111)
||(x_pointer == 54 && y_pointer == 111)
||(x_pointer == 55 && y_pointer == 111)
||(x_pointer == 56 && y_pointer == 111)
||(x_pointer == 57 && y_pointer == 111)
||(x_pointer == 58 && y_pointer == 111)
||(x_pointer == 59 && y_pointer == 111)
||(x_pointer == 60 && y_pointer == 111)
||(x_pointer == 61 && y_pointer == 111)
||(x_pointer == 62 && y_pointer == 111)
||(x_pointer == 63 && y_pointer == 111)
||(x_pointer == 64 && y_pointer == 111)
||(x_pointer == 65 && y_pointer == 111)
||(x_pointer == 66 && y_pointer == 111)
||(x_pointer == 67 && y_pointer == 111)
||(x_pointer == 68 && y_pointer == 111)
||(x_pointer == 69 && y_pointer == 111)
||(x_pointer == 70 && y_pointer == 111)
||(x_pointer == 71 && y_pointer == 111)
||(x_pointer == 72 && y_pointer == 111)
||(x_pointer == 73 && y_pointer == 111)
||(x_pointer == 74 && y_pointer == 111)
||(x_pointer == 75 && y_pointer == 111)
||(x_pointer == 76 && y_pointer == 111)
||(x_pointer == 77 && y_pointer == 111)
||(x_pointer == 78 && y_pointer == 111)
||(x_pointer == 79 && y_pointer == 111)
||(x_pointer == 80 && y_pointer == 111)
||(x_pointer == 81 && y_pointer == 111)
||(x_pointer == 82 && y_pointer == 111)
||(x_pointer == 83 && y_pointer == 111)
||(x_pointer == 84 && y_pointer == 111)
||(x_pointer == 85 && y_pointer == 111)
||(x_pointer == 86 && y_pointer == 111)
||(x_pointer == 87 && y_pointer == 111)
||(x_pointer == 88 && y_pointer == 111)
||(x_pointer == 89 && y_pointer == 111)
||(x_pointer == 90 && y_pointer == 111)
||(x_pointer == 91 && y_pointer == 111)
||(x_pointer == 92 && y_pointer == 111)
||(x_pointer == 93 && y_pointer == 111)
||(x_pointer == 94 && y_pointer == 111)
||(x_pointer == 95 && y_pointer == 111)
||(x_pointer == 96 && y_pointer == 111)
||(x_pointer == 97 && y_pointer == 111)
||(x_pointer == 98 && y_pointer == 111)
||(x_pointer == 99 && y_pointer == 111)
||(x_pointer == 100 && y_pointer == 111)
||(x_pointer == 101 && y_pointer == 111)
||(x_pointer == 102 && y_pointer == 111)
||(x_pointer == 103 && y_pointer == 111)
||(x_pointer == 104 && y_pointer == 111)
||(x_pointer == 105 && y_pointer == 111)
||(x_pointer == 106 && y_pointer == 111)
||(x_pointer == 107 && y_pointer == 111)
||(x_pointer == 108 && y_pointer == 111)
||(x_pointer == 109 && y_pointer == 111)
||(x_pointer == 110 && y_pointer == 111)
||(x_pointer == 111 && y_pointer == 111)
||(x_pointer == 112 && y_pointer == 111)
||(x_pointer == 113 && y_pointer == 111)
||(x_pointer == 114 && y_pointer == 111)
||(x_pointer == 115 && y_pointer == 111)
||(x_pointer == 116 && y_pointer == 111)
||(x_pointer == 117 && y_pointer == 111)
||(x_pointer == 118 && y_pointer == 111)
||(x_pointer == 119 && y_pointer == 111)
||(x_pointer == 120 && y_pointer == 111)
||(x_pointer == 121 && y_pointer == 111)
||(x_pointer == 122 && y_pointer == 111)
||(x_pointer == 123 && y_pointer == 111)
||(x_pointer == 124 && y_pointer == 111)
||(x_pointer == 125 && y_pointer == 111)
||(x_pointer == 126 && y_pointer == 111)
||(x_pointer == 127 && y_pointer == 111)
||(x_pointer == 128 && y_pointer == 111)
||(x_pointer == 129 && y_pointer == 111)
||(x_pointer == 130 && y_pointer == 111)
||(x_pointer == 131 && y_pointer == 111)
||(x_pointer == 132 && y_pointer == 111)
||(x_pointer == 133 && y_pointer == 111)
||(x_pointer == 134 && y_pointer == 111)
||(x_pointer == 135 && y_pointer == 111)
||(x_pointer == 136 && y_pointer == 111)
||(x_pointer == 137 && y_pointer == 111)
||(x_pointer == 138 && y_pointer == 111)
||(x_pointer == 139 && y_pointer == 111)
||(x_pointer == 140 && y_pointer == 111)
||(x_pointer == 141 && y_pointer == 111)
||(x_pointer == 142 && y_pointer == 111)
||(x_pointer == 143 && y_pointer == 111)
||(x_pointer == 144 && y_pointer == 111)
||(x_pointer == 145 && y_pointer == 111)
||(x_pointer == 146 && y_pointer == 111)
||(x_pointer == 147 && y_pointer == 111)
||(x_pointer == 148 && y_pointer == 111)
||(x_pointer == 149 && y_pointer == 111)
||(x_pointer == 150 && y_pointer == 111)
||(x_pointer == 151 && y_pointer == 111)
||(x_pointer == 152 && y_pointer == 111)
||(x_pointer == 153 && y_pointer == 111)
||(x_pointer == 154 && y_pointer == 111)
||(x_pointer == 155 && y_pointer == 111)
||(x_pointer == 156 && y_pointer == 111)
||(x_pointer == 157 && y_pointer == 111)
||(x_pointer == 2 && y_pointer == 112)
||(x_pointer == 3 && y_pointer == 112)
||(x_pointer == 4 && y_pointer == 112)
||(x_pointer == 5 && y_pointer == 112)
||(x_pointer == 6 && y_pointer == 112)
||(x_pointer == 7 && y_pointer == 112)
||(x_pointer == 8 && y_pointer == 112)
||(x_pointer == 9 && y_pointer == 112)
||(x_pointer == 10 && y_pointer == 112)
||(x_pointer == 11 && y_pointer == 112)
||(x_pointer == 12 && y_pointer == 112)
||(x_pointer == 13 && y_pointer == 112)
||(x_pointer == 14 && y_pointer == 112)
||(x_pointer == 15 && y_pointer == 112)
||(x_pointer == 16 && y_pointer == 112)
||(x_pointer == 17 && y_pointer == 112)
||(x_pointer == 18 && y_pointer == 112)
||(x_pointer == 19 && y_pointer == 112)
||(x_pointer == 20 && y_pointer == 112)
||(x_pointer == 21 && y_pointer == 112)
||(x_pointer == 22 && y_pointer == 112)
||(x_pointer == 23 && y_pointer == 112)
||(x_pointer == 24 && y_pointer == 112)
||(x_pointer == 25 && y_pointer == 112)
||(x_pointer == 26 && y_pointer == 112)
||(x_pointer == 27 && y_pointer == 112)
||(x_pointer == 28 && y_pointer == 112)
||(x_pointer == 29 && y_pointer == 112)
||(x_pointer == 30 && y_pointer == 112)
||(x_pointer == 31 && y_pointer == 112)
||(x_pointer == 32 && y_pointer == 112)
||(x_pointer == 33 && y_pointer == 112)
||(x_pointer == 34 && y_pointer == 112)
||(x_pointer == 35 && y_pointer == 112)
||(x_pointer == 36 && y_pointer == 112)
||(x_pointer == 37 && y_pointer == 112)
||(x_pointer == 38 && y_pointer == 112)
||(x_pointer == 39 && y_pointer == 112)
||(x_pointer == 40 && y_pointer == 112)
||(x_pointer == 41 && y_pointer == 112)
||(x_pointer == 42 && y_pointer == 112)
||(x_pointer == 43 && y_pointer == 112)
||(x_pointer == 44 && y_pointer == 112)
||(x_pointer == 45 && y_pointer == 112)
||(x_pointer == 46 && y_pointer == 112)
||(x_pointer == 47 && y_pointer == 112)
||(x_pointer == 48 && y_pointer == 112)
||(x_pointer == 49 && y_pointer == 112)
||(x_pointer == 50 && y_pointer == 112)
||(x_pointer == 51 && y_pointer == 112)
||(x_pointer == 52 && y_pointer == 112)
||(x_pointer == 53 && y_pointer == 112)
||(x_pointer == 54 && y_pointer == 112)
||(x_pointer == 55 && y_pointer == 112)
||(x_pointer == 56 && y_pointer == 112)
||(x_pointer == 57 && y_pointer == 112)
||(x_pointer == 58 && y_pointer == 112)
||(x_pointer == 59 && y_pointer == 112)
||(x_pointer == 60 && y_pointer == 112)
||(x_pointer == 61 && y_pointer == 112)
||(x_pointer == 62 && y_pointer == 112)
||(x_pointer == 63 && y_pointer == 112)
||(x_pointer == 64 && y_pointer == 112)
||(x_pointer == 65 && y_pointer == 112)
||(x_pointer == 66 && y_pointer == 112)
||(x_pointer == 67 && y_pointer == 112)
||(x_pointer == 68 && y_pointer == 112)
||(x_pointer == 69 && y_pointer == 112)
||(x_pointer == 70 && y_pointer == 112)
||(x_pointer == 71 && y_pointer == 112)
||(x_pointer == 72 && y_pointer == 112)
||(x_pointer == 73 && y_pointer == 112)
||(x_pointer == 74 && y_pointer == 112)
||(x_pointer == 75 && y_pointer == 112)
||(x_pointer == 76 && y_pointer == 112)
||(x_pointer == 77 && y_pointer == 112)
||(x_pointer == 78 && y_pointer == 112)
||(x_pointer == 79 && y_pointer == 112)
||(x_pointer == 80 && y_pointer == 112)
||(x_pointer == 81 && y_pointer == 112)
||(x_pointer == 82 && y_pointer == 112)
||(x_pointer == 83 && y_pointer == 112)
||(x_pointer == 84 && y_pointer == 112)
||(x_pointer == 85 && y_pointer == 112)
||(x_pointer == 86 && y_pointer == 112)
||(x_pointer == 87 && y_pointer == 112)
||(x_pointer == 88 && y_pointer == 112)
||(x_pointer == 89 && y_pointer == 112)
||(x_pointer == 90 && y_pointer == 112)
||(x_pointer == 91 && y_pointer == 112)
||(x_pointer == 92 && y_pointer == 112)
||(x_pointer == 93 && y_pointer == 112)
||(x_pointer == 94 && y_pointer == 112)
||(x_pointer == 95 && y_pointer == 112)
||(x_pointer == 96 && y_pointer == 112)
||(x_pointer == 97 && y_pointer == 112)
||(x_pointer == 98 && y_pointer == 112)
||(x_pointer == 99 && y_pointer == 112)
||(x_pointer == 100 && y_pointer == 112)
||(x_pointer == 101 && y_pointer == 112)
||(x_pointer == 102 && y_pointer == 112)
||(x_pointer == 103 && y_pointer == 112)
||(x_pointer == 104 && y_pointer == 112)
||(x_pointer == 105 && y_pointer == 112)
||(x_pointer == 106 && y_pointer == 112)
||(x_pointer == 107 && y_pointer == 112)
||(x_pointer == 108 && y_pointer == 112)
||(x_pointer == 109 && y_pointer == 112)
||(x_pointer == 110 && y_pointer == 112)
||(x_pointer == 111 && y_pointer == 112)
||(x_pointer == 112 && y_pointer == 112)
||(x_pointer == 113 && y_pointer == 112)
||(x_pointer == 114 && y_pointer == 112)
||(x_pointer == 115 && y_pointer == 112)
||(x_pointer == 116 && y_pointer == 112)
||(x_pointer == 117 && y_pointer == 112)
||(x_pointer == 118 && y_pointer == 112)
||(x_pointer == 119 && y_pointer == 112)
||(x_pointer == 120 && y_pointer == 112)
||(x_pointer == 121 && y_pointer == 112)
||(x_pointer == 122 && y_pointer == 112)
||(x_pointer == 123 && y_pointer == 112)
||(x_pointer == 124 && y_pointer == 112)
||(x_pointer == 125 && y_pointer == 112)
||(x_pointer == 126 && y_pointer == 112)
||(x_pointer == 127 && y_pointer == 112)
||(x_pointer == 128 && y_pointer == 112)
||(x_pointer == 129 && y_pointer == 112)
||(x_pointer == 130 && y_pointer == 112)
||(x_pointer == 131 && y_pointer == 112)
||(x_pointer == 132 && y_pointer == 112)
||(x_pointer == 133 && y_pointer == 112)
||(x_pointer == 134 && y_pointer == 112)
||(x_pointer == 135 && y_pointer == 112)
||(x_pointer == 136 && y_pointer == 112)
||(x_pointer == 137 && y_pointer == 112)
||(x_pointer == 138 && y_pointer == 112)
||(x_pointer == 139 && y_pointer == 112)
||(x_pointer == 140 && y_pointer == 112)
||(x_pointer == 141 && y_pointer == 112)
||(x_pointer == 142 && y_pointer == 112)
||(x_pointer == 143 && y_pointer == 112)
||(x_pointer == 144 && y_pointer == 112)
||(x_pointer == 145 && y_pointer == 112)
||(x_pointer == 146 && y_pointer == 112)
||(x_pointer == 147 && y_pointer == 112)
||(x_pointer == 148 && y_pointer == 112)
||(x_pointer == 149 && y_pointer == 112)
||(x_pointer == 150 && y_pointer == 112)
||(x_pointer == 151 && y_pointer == 112)
||(x_pointer == 152 && y_pointer == 112)
||(x_pointer == 153 && y_pointer == 112)
||(x_pointer == 154 && y_pointer == 112)
||(x_pointer == 155 && y_pointer == 112)
||(x_pointer == 156 && y_pointer == 112)
||(x_pointer == 157 && y_pointer == 112));
	
	wire barrier_pixel_3 = current_level == 3 && ((x_pointer == 23 && y_pointer == 14)
||(x_pointer == 24 && y_pointer == 14)
||(x_pointer == 25 && y_pointer == 14)
||(x_pointer == 26 && y_pointer == 14)
||(x_pointer == 27 && y_pointer == 14)
||(x_pointer == 28 && y_pointer == 14)
||(x_pointer == 29 && y_pointer == 14)
||(x_pointer == 30 && y_pointer == 14)
||(x_pointer == 31 && y_pointer == 14)
||(x_pointer == 32 && y_pointer == 14)
||(x_pointer == 33 && y_pointer == 14)
||(x_pointer == 34 && y_pointer == 14)
||(x_pointer == 35 && y_pointer == 14)
||(x_pointer == 36 && y_pointer == 14)
||(x_pointer == 37 && y_pointer == 14)
||(x_pointer == 38 && y_pointer == 14)
||(x_pointer == 39 && y_pointer == 14)
||(x_pointer == 40 && y_pointer == 14)
||(x_pointer == 41 && y_pointer == 14)
||(x_pointer == 42 && y_pointer == 14)
||(x_pointer == 43 && y_pointer == 14)
||(x_pointer == 122 && y_pointer == 14)
||(x_pointer == 123 && y_pointer == 14)
||(x_pointer == 124 && y_pointer == 14)
||(x_pointer == 125 && y_pointer == 14)
||(x_pointer == 126 && y_pointer == 14)
||(x_pointer == 127 && y_pointer == 14)
||(x_pointer == 128 && y_pointer == 14)
||(x_pointer == 129 && y_pointer == 14)
||(x_pointer == 130 && y_pointer == 14)
||(x_pointer == 131 && y_pointer == 14)
||(x_pointer == 132 && y_pointer == 14)
||(x_pointer == 133 && y_pointer == 14)
||(x_pointer == 134 && y_pointer == 14)
||(x_pointer == 135 && y_pointer == 14)
||(x_pointer == 136 && y_pointer == 14)
||(x_pointer == 137 && y_pointer == 14)
||(x_pointer == 138 && y_pointer == 14)
||(x_pointer == 139 && y_pointer == 14)
||(x_pointer == 140 && y_pointer == 14)
||(x_pointer == 141 && y_pointer == 14)
||(x_pointer == 142 && y_pointer == 14)
||(x_pointer == 23 && y_pointer == 15)
||(x_pointer == 24 && y_pointer == 15)
||(x_pointer == 25 && y_pointer == 15)
||(x_pointer == 26 && y_pointer == 15)
||(x_pointer == 27 && y_pointer == 15)
||(x_pointer == 28 && y_pointer == 15)
||(x_pointer == 29 && y_pointer == 15)
||(x_pointer == 30 && y_pointer == 15)
||(x_pointer == 31 && y_pointer == 15)
||(x_pointer == 32 && y_pointer == 15)
||(x_pointer == 33 && y_pointer == 15)
||(x_pointer == 34 && y_pointer == 15)
||(x_pointer == 35 && y_pointer == 15)
||(x_pointer == 36 && y_pointer == 15)
||(x_pointer == 37 && y_pointer == 15)
||(x_pointer == 38 && y_pointer == 15)
||(x_pointer == 39 && y_pointer == 15)
||(x_pointer == 40 && y_pointer == 15)
||(x_pointer == 41 && y_pointer == 15)
||(x_pointer == 42 && y_pointer == 15)
||(x_pointer == 43 && y_pointer == 15)
||(x_pointer == 122 && y_pointer == 15)
||(x_pointer == 123 && y_pointer == 15)
||(x_pointer == 124 && y_pointer == 15)
||(x_pointer == 125 && y_pointer == 15)
||(x_pointer == 126 && y_pointer == 15)
||(x_pointer == 127 && y_pointer == 15)
||(x_pointer == 128 && y_pointer == 15)
||(x_pointer == 129 && y_pointer == 15)
||(x_pointer == 130 && y_pointer == 15)
||(x_pointer == 131 && y_pointer == 15)
||(x_pointer == 132 && y_pointer == 15)
||(x_pointer == 133 && y_pointer == 15)
||(x_pointer == 134 && y_pointer == 15)
||(x_pointer == 135 && y_pointer == 15)
||(x_pointer == 136 && y_pointer == 15)
||(x_pointer == 137 && y_pointer == 15)
||(x_pointer == 138 && y_pointer == 15)
||(x_pointer == 139 && y_pointer == 15)
||(x_pointer == 140 && y_pointer == 15)
||(x_pointer == 141 && y_pointer == 15)
||(x_pointer == 142 && y_pointer == 15)
||(x_pointer == 23 && y_pointer == 16)
||(x_pointer == 24 && y_pointer == 16)
||(x_pointer == 25 && y_pointer == 16)
||(x_pointer == 26 && y_pointer == 16)
||(x_pointer == 27 && y_pointer == 16)
||(x_pointer == 28 && y_pointer == 16)
||(x_pointer == 29 && y_pointer == 16)
||(x_pointer == 30 && y_pointer == 16)
||(x_pointer == 31 && y_pointer == 16)
||(x_pointer == 32 && y_pointer == 16)
||(x_pointer == 33 && y_pointer == 16)
||(x_pointer == 34 && y_pointer == 16)
||(x_pointer == 35 && y_pointer == 16)
||(x_pointer == 36 && y_pointer == 16)
||(x_pointer == 37 && y_pointer == 16)
||(x_pointer == 38 && y_pointer == 16)
||(x_pointer == 39 && y_pointer == 16)
||(x_pointer == 40 && y_pointer == 16)
||(x_pointer == 41 && y_pointer == 16)
||(x_pointer == 42 && y_pointer == 16)
||(x_pointer == 43 && y_pointer == 16)
||(x_pointer == 122 && y_pointer == 16)
||(x_pointer == 123 && y_pointer == 16)
||(x_pointer == 124 && y_pointer == 16)
||(x_pointer == 125 && y_pointer == 16)
||(x_pointer == 126 && y_pointer == 16)
||(x_pointer == 127 && y_pointer == 16)
||(x_pointer == 128 && y_pointer == 16)
||(x_pointer == 129 && y_pointer == 16)
||(x_pointer == 130 && y_pointer == 16)
||(x_pointer == 131 && y_pointer == 16)
||(x_pointer == 132 && y_pointer == 16)
||(x_pointer == 133 && y_pointer == 16)
||(x_pointer == 134 && y_pointer == 16)
||(x_pointer == 135 && y_pointer == 16)
||(x_pointer == 136 && y_pointer == 16)
||(x_pointer == 137 && y_pointer == 16)
||(x_pointer == 138 && y_pointer == 16)
||(x_pointer == 139 && y_pointer == 16)
||(x_pointer == 140 && y_pointer == 16)
||(x_pointer == 141 && y_pointer == 16)
||(x_pointer == 142 && y_pointer == 16)
||(x_pointer == 23 && y_pointer == 17)
||(x_pointer == 24 && y_pointer == 17)
||(x_pointer == 25 && y_pointer == 17)
||(x_pointer == 26 && y_pointer == 17)
||(x_pointer == 27 && y_pointer == 17)
||(x_pointer == 28 && y_pointer == 17)
||(x_pointer == 29 && y_pointer == 17)
||(x_pointer == 30 && y_pointer == 17)
||(x_pointer == 31 && y_pointer == 17)
||(x_pointer == 32 && y_pointer == 17)
||(x_pointer == 33 && y_pointer == 17)
||(x_pointer == 34 && y_pointer == 17)
||(x_pointer == 35 && y_pointer == 17)
||(x_pointer == 36 && y_pointer == 17)
||(x_pointer == 37 && y_pointer == 17)
||(x_pointer == 38 && y_pointer == 17)
||(x_pointer == 39 && y_pointer == 17)
||(x_pointer == 40 && y_pointer == 17)
||(x_pointer == 41 && y_pointer == 17)
||(x_pointer == 42 && y_pointer == 17)
||(x_pointer == 43 && y_pointer == 17)
||(x_pointer == 122 && y_pointer == 17)
||(x_pointer == 123 && y_pointer == 17)
||(x_pointer == 124 && y_pointer == 17)
||(x_pointer == 125 && y_pointer == 17)
||(x_pointer == 126 && y_pointer == 17)
||(x_pointer == 127 && y_pointer == 17)
||(x_pointer == 128 && y_pointer == 17)
||(x_pointer == 129 && y_pointer == 17)
||(x_pointer == 130 && y_pointer == 17)
||(x_pointer == 131 && y_pointer == 17)
||(x_pointer == 132 && y_pointer == 17)
||(x_pointer == 133 && y_pointer == 17)
||(x_pointer == 134 && y_pointer == 17)
||(x_pointer == 135 && y_pointer == 17)
||(x_pointer == 136 && y_pointer == 17)
||(x_pointer == 137 && y_pointer == 17)
||(x_pointer == 138 && y_pointer == 17)
||(x_pointer == 139 && y_pointer == 17)
||(x_pointer == 140 && y_pointer == 17)
||(x_pointer == 141 && y_pointer == 17)
||(x_pointer == 142 && y_pointer == 17)
||(x_pointer == 23 && y_pointer == 18)
||(x_pointer == 24 && y_pointer == 18)
||(x_pointer == 25 && y_pointer == 18)
||(x_pointer == 26 && y_pointer == 18)
||(x_pointer == 27 && y_pointer == 18)
||(x_pointer == 28 && y_pointer == 18)
||(x_pointer == 29 && y_pointer == 18)
||(x_pointer == 30 && y_pointer == 18)
||(x_pointer == 31 && y_pointer == 18)
||(x_pointer == 32 && y_pointer == 18)
||(x_pointer == 33 && y_pointer == 18)
||(x_pointer == 34 && y_pointer == 18)
||(x_pointer == 35 && y_pointer == 18)
||(x_pointer == 36 && y_pointer == 18)
||(x_pointer == 37 && y_pointer == 18)
||(x_pointer == 38 && y_pointer == 18)
||(x_pointer == 39 && y_pointer == 18)
||(x_pointer == 40 && y_pointer == 18)
||(x_pointer == 41 && y_pointer == 18)
||(x_pointer == 42 && y_pointer == 18)
||(x_pointer == 43 && y_pointer == 18)
||(x_pointer == 122 && y_pointer == 18)
||(x_pointer == 123 && y_pointer == 18)
||(x_pointer == 124 && y_pointer == 18)
||(x_pointer == 125 && y_pointer == 18)
||(x_pointer == 126 && y_pointer == 18)
||(x_pointer == 127 && y_pointer == 18)
||(x_pointer == 128 && y_pointer == 18)
||(x_pointer == 129 && y_pointer == 18)
||(x_pointer == 130 && y_pointer == 18)
||(x_pointer == 131 && y_pointer == 18)
||(x_pointer == 132 && y_pointer == 18)
||(x_pointer == 133 && y_pointer == 18)
||(x_pointer == 134 && y_pointer == 18)
||(x_pointer == 135 && y_pointer == 18)
||(x_pointer == 136 && y_pointer == 18)
||(x_pointer == 137 && y_pointer == 18)
||(x_pointer == 138 && y_pointer == 18)
||(x_pointer == 139 && y_pointer == 18)
||(x_pointer == 140 && y_pointer == 18)
||(x_pointer == 141 && y_pointer == 18)
||(x_pointer == 142 && y_pointer == 18)
||(x_pointer == 23 && y_pointer == 19)
||(x_pointer == 24 && y_pointer == 19)
||(x_pointer == 25 && y_pointer == 19)
||(x_pointer == 26 && y_pointer == 19)
||(x_pointer == 27 && y_pointer == 19)
||(x_pointer == 28 && y_pointer == 19)
||(x_pointer == 29 && y_pointer == 19)
||(x_pointer == 30 && y_pointer == 19)
||(x_pointer == 31 && y_pointer == 19)
||(x_pointer == 32 && y_pointer == 19)
||(x_pointer == 33 && y_pointer == 19)
||(x_pointer == 34 && y_pointer == 19)
||(x_pointer == 35 && y_pointer == 19)
||(x_pointer == 36 && y_pointer == 19)
||(x_pointer == 37 && y_pointer == 19)
||(x_pointer == 38 && y_pointer == 19)
||(x_pointer == 39 && y_pointer == 19)
||(x_pointer == 40 && y_pointer == 19)
||(x_pointer == 41 && y_pointer == 19)
||(x_pointer == 42 && y_pointer == 19)
||(x_pointer == 43 && y_pointer == 19)
||(x_pointer == 122 && y_pointer == 19)
||(x_pointer == 123 && y_pointer == 19)
||(x_pointer == 124 && y_pointer == 19)
||(x_pointer == 125 && y_pointer == 19)
||(x_pointer == 126 && y_pointer == 19)
||(x_pointer == 127 && y_pointer == 19)
||(x_pointer == 128 && y_pointer == 19)
||(x_pointer == 129 && y_pointer == 19)
||(x_pointer == 130 && y_pointer == 19)
||(x_pointer == 131 && y_pointer == 19)
||(x_pointer == 132 && y_pointer == 19)
||(x_pointer == 133 && y_pointer == 19)
||(x_pointer == 134 && y_pointer == 19)
||(x_pointer == 135 && y_pointer == 19)
||(x_pointer == 136 && y_pointer == 19)
||(x_pointer == 137 && y_pointer == 19)
||(x_pointer == 138 && y_pointer == 19)
||(x_pointer == 139 && y_pointer == 19)
||(x_pointer == 140 && y_pointer == 19)
||(x_pointer == 141 && y_pointer == 19)
||(x_pointer == 142 && y_pointer == 19)
||(x_pointer == 23 && y_pointer == 20)
||(x_pointer == 24 && y_pointer == 20)
||(x_pointer == 25 && y_pointer == 20)
||(x_pointer == 26 && y_pointer == 20)
||(x_pointer == 27 && y_pointer == 20)
||(x_pointer == 28 && y_pointer == 20)
||(x_pointer == 29 && y_pointer == 20)
||(x_pointer == 30 && y_pointer == 20)
||(x_pointer == 31 && y_pointer == 20)
||(x_pointer == 32 && y_pointer == 20)
||(x_pointer == 33 && y_pointer == 20)
||(x_pointer == 34 && y_pointer == 20)
||(x_pointer == 35 && y_pointer == 20)
||(x_pointer == 36 && y_pointer == 20)
||(x_pointer == 37 && y_pointer == 20)
||(x_pointer == 38 && y_pointer == 20)
||(x_pointer == 39 && y_pointer == 20)
||(x_pointer == 40 && y_pointer == 20)
||(x_pointer == 41 && y_pointer == 20)
||(x_pointer == 42 && y_pointer == 20)
||(x_pointer == 43 && y_pointer == 20)
||(x_pointer == 122 && y_pointer == 20)
||(x_pointer == 123 && y_pointer == 20)
||(x_pointer == 124 && y_pointer == 20)
||(x_pointer == 125 && y_pointer == 20)
||(x_pointer == 126 && y_pointer == 20)
||(x_pointer == 127 && y_pointer == 20)
||(x_pointer == 128 && y_pointer == 20)
||(x_pointer == 129 && y_pointer == 20)
||(x_pointer == 130 && y_pointer == 20)
||(x_pointer == 131 && y_pointer == 20)
||(x_pointer == 132 && y_pointer == 20)
||(x_pointer == 133 && y_pointer == 20)
||(x_pointer == 134 && y_pointer == 20)
||(x_pointer == 135 && y_pointer == 20)
||(x_pointer == 136 && y_pointer == 20)
||(x_pointer == 137 && y_pointer == 20)
||(x_pointer == 138 && y_pointer == 20)
||(x_pointer == 139 && y_pointer == 20)
||(x_pointer == 140 && y_pointer == 20)
||(x_pointer == 141 && y_pointer == 20)
||(x_pointer == 142 && y_pointer == 20)
||(x_pointer == 23 && y_pointer == 21)
||(x_pointer == 24 && y_pointer == 21)
||(x_pointer == 25 && y_pointer == 21)
||(x_pointer == 26 && y_pointer == 21)
||(x_pointer == 27 && y_pointer == 21)
||(x_pointer == 28 && y_pointer == 21)
||(x_pointer == 29 && y_pointer == 21)
||(x_pointer == 30 && y_pointer == 21)
||(x_pointer == 31 && y_pointer == 21)
||(x_pointer == 32 && y_pointer == 21)
||(x_pointer == 33 && y_pointer == 21)
||(x_pointer == 34 && y_pointer == 21)
||(x_pointer == 35 && y_pointer == 21)
||(x_pointer == 36 && y_pointer == 21)
||(x_pointer == 37 && y_pointer == 21)
||(x_pointer == 38 && y_pointer == 21)
||(x_pointer == 39 && y_pointer == 21)
||(x_pointer == 40 && y_pointer == 21)
||(x_pointer == 41 && y_pointer == 21)
||(x_pointer == 42 && y_pointer == 21)
||(x_pointer == 43 && y_pointer == 21)
||(x_pointer == 122 && y_pointer == 21)
||(x_pointer == 123 && y_pointer == 21)
||(x_pointer == 124 && y_pointer == 21)
||(x_pointer == 125 && y_pointer == 21)
||(x_pointer == 126 && y_pointer == 21)
||(x_pointer == 127 && y_pointer == 21)
||(x_pointer == 128 && y_pointer == 21)
||(x_pointer == 129 && y_pointer == 21)
||(x_pointer == 130 && y_pointer == 21)
||(x_pointer == 131 && y_pointer == 21)
||(x_pointer == 132 && y_pointer == 21)
||(x_pointer == 133 && y_pointer == 21)
||(x_pointer == 134 && y_pointer == 21)
||(x_pointer == 135 && y_pointer == 21)
||(x_pointer == 136 && y_pointer == 21)
||(x_pointer == 137 && y_pointer == 21)
||(x_pointer == 138 && y_pointer == 21)
||(x_pointer == 139 && y_pointer == 21)
||(x_pointer == 140 && y_pointer == 21)
||(x_pointer == 141 && y_pointer == 21)
||(x_pointer == 142 && y_pointer == 21)
||(x_pointer == 23 && y_pointer == 22)
||(x_pointer == 24 && y_pointer == 22)
||(x_pointer == 25 && y_pointer == 22)
||(x_pointer == 26 && y_pointer == 22)
||(x_pointer == 27 && y_pointer == 22)
||(x_pointer == 28 && y_pointer == 22)
||(x_pointer == 29 && y_pointer == 22)
||(x_pointer == 30 && y_pointer == 22)
||(x_pointer == 31 && y_pointer == 22)
||(x_pointer == 32 && y_pointer == 22)
||(x_pointer == 33 && y_pointer == 22)
||(x_pointer == 34 && y_pointer == 22)
||(x_pointer == 35 && y_pointer == 22)
||(x_pointer == 36 && y_pointer == 22)
||(x_pointer == 37 && y_pointer == 22)
||(x_pointer == 38 && y_pointer == 22)
||(x_pointer == 39 && y_pointer == 22)
||(x_pointer == 40 && y_pointer == 22)
||(x_pointer == 41 && y_pointer == 22)
||(x_pointer == 42 && y_pointer == 22)
||(x_pointer == 43 && y_pointer == 22)
||(x_pointer == 122 && y_pointer == 22)
||(x_pointer == 123 && y_pointer == 22)
||(x_pointer == 124 && y_pointer == 22)
||(x_pointer == 125 && y_pointer == 22)
||(x_pointer == 126 && y_pointer == 22)
||(x_pointer == 127 && y_pointer == 22)
||(x_pointer == 128 && y_pointer == 22)
||(x_pointer == 129 && y_pointer == 22)
||(x_pointer == 130 && y_pointer == 22)
||(x_pointer == 131 && y_pointer == 22)
||(x_pointer == 132 && y_pointer == 22)
||(x_pointer == 133 && y_pointer == 22)
||(x_pointer == 134 && y_pointer == 22)
||(x_pointer == 135 && y_pointer == 22)
||(x_pointer == 136 && y_pointer == 22)
||(x_pointer == 137 && y_pointer == 22)
||(x_pointer == 138 && y_pointer == 22)
||(x_pointer == 139 && y_pointer == 22)
||(x_pointer == 140 && y_pointer == 22)
||(x_pointer == 141 && y_pointer == 22)
||(x_pointer == 142 && y_pointer == 22)
||(x_pointer == 23 && y_pointer == 23)
||(x_pointer == 24 && y_pointer == 23)
||(x_pointer == 25 && y_pointer == 23)
||(x_pointer == 26 && y_pointer == 23)
||(x_pointer == 27 && y_pointer == 23)
||(x_pointer == 28 && y_pointer == 23)
||(x_pointer == 29 && y_pointer == 23)
||(x_pointer == 30 && y_pointer == 23)
||(x_pointer == 31 && y_pointer == 23)
||(x_pointer == 134 && y_pointer == 23)
||(x_pointer == 135 && y_pointer == 23)
||(x_pointer == 136 && y_pointer == 23)
||(x_pointer == 137 && y_pointer == 23)
||(x_pointer == 138 && y_pointer == 23)
||(x_pointer == 139 && y_pointer == 23)
||(x_pointer == 140 && y_pointer == 23)
||(x_pointer == 141 && y_pointer == 23)
||(x_pointer == 142 && y_pointer == 23)
||(x_pointer == 23 && y_pointer == 24)
||(x_pointer == 24 && y_pointer == 24)
||(x_pointer == 25 && y_pointer == 24)
||(x_pointer == 26 && y_pointer == 24)
||(x_pointer == 27 && y_pointer == 24)
||(x_pointer == 28 && y_pointer == 24)
||(x_pointer == 29 && y_pointer == 24)
||(x_pointer == 30 && y_pointer == 24)
||(x_pointer == 31 && y_pointer == 24)
||(x_pointer == 134 && y_pointer == 24)
||(x_pointer == 135 && y_pointer == 24)
||(x_pointer == 136 && y_pointer == 24)
||(x_pointer == 137 && y_pointer == 24)
||(x_pointer == 138 && y_pointer == 24)
||(x_pointer == 139 && y_pointer == 24)
||(x_pointer == 140 && y_pointer == 24)
||(x_pointer == 141 && y_pointer == 24)
||(x_pointer == 142 && y_pointer == 24)
||(x_pointer == 23 && y_pointer == 25)
||(x_pointer == 24 && y_pointer == 25)
||(x_pointer == 25 && y_pointer == 25)
||(x_pointer == 26 && y_pointer == 25)
||(x_pointer == 27 && y_pointer == 25)
||(x_pointer == 28 && y_pointer == 25)
||(x_pointer == 29 && y_pointer == 25)
||(x_pointer == 30 && y_pointer == 25)
||(x_pointer == 31 && y_pointer == 25)
||(x_pointer == 134 && y_pointer == 25)
||(x_pointer == 135 && y_pointer == 25)
||(x_pointer == 136 && y_pointer == 25)
||(x_pointer == 137 && y_pointer == 25)
||(x_pointer == 138 && y_pointer == 25)
||(x_pointer == 139 && y_pointer == 25)
||(x_pointer == 140 && y_pointer == 25)
||(x_pointer == 141 && y_pointer == 25)
||(x_pointer == 142 && y_pointer == 25)
||(x_pointer == 23 && y_pointer == 26)
||(x_pointer == 24 && y_pointer == 26)
||(x_pointer == 25 && y_pointer == 26)
||(x_pointer == 26 && y_pointer == 26)
||(x_pointer == 27 && y_pointer == 26)
||(x_pointer == 28 && y_pointer == 26)
||(x_pointer == 29 && y_pointer == 26)
||(x_pointer == 30 && y_pointer == 26)
||(x_pointer == 31 && y_pointer == 26)
||(x_pointer == 134 && y_pointer == 26)
||(x_pointer == 135 && y_pointer == 26)
||(x_pointer == 136 && y_pointer == 26)
||(x_pointer == 137 && y_pointer == 26)
||(x_pointer == 138 && y_pointer == 26)
||(x_pointer == 139 && y_pointer == 26)
||(x_pointer == 140 && y_pointer == 26)
||(x_pointer == 141 && y_pointer == 26)
||(x_pointer == 142 && y_pointer == 26)
||(x_pointer == 23 && y_pointer == 27)
||(x_pointer == 24 && y_pointer == 27)
||(x_pointer == 25 && y_pointer == 27)
||(x_pointer == 26 && y_pointer == 27)
||(x_pointer == 27 && y_pointer == 27)
||(x_pointer == 28 && y_pointer == 27)
||(x_pointer == 29 && y_pointer == 27)
||(x_pointer == 30 && y_pointer == 27)
||(x_pointer == 31 && y_pointer == 27)
||(x_pointer == 134 && y_pointer == 27)
||(x_pointer == 135 && y_pointer == 27)
||(x_pointer == 136 && y_pointer == 27)
||(x_pointer == 137 && y_pointer == 27)
||(x_pointer == 138 && y_pointer == 27)
||(x_pointer == 139 && y_pointer == 27)
||(x_pointer == 140 && y_pointer == 27)
||(x_pointer == 141 && y_pointer == 27)
||(x_pointer == 142 && y_pointer == 27)
||(x_pointer == 23 && y_pointer == 28)
||(x_pointer == 24 && y_pointer == 28)
||(x_pointer == 25 && y_pointer == 28)
||(x_pointer == 26 && y_pointer == 28)
||(x_pointer == 27 && y_pointer == 28)
||(x_pointer == 28 && y_pointer == 28)
||(x_pointer == 29 && y_pointer == 28)
||(x_pointer == 30 && y_pointer == 28)
||(x_pointer == 31 && y_pointer == 28)
||(x_pointer == 134 && y_pointer == 28)
||(x_pointer == 135 && y_pointer == 28)
||(x_pointer == 136 && y_pointer == 28)
||(x_pointer == 137 && y_pointer == 28)
||(x_pointer == 138 && y_pointer == 28)
||(x_pointer == 139 && y_pointer == 28)
||(x_pointer == 140 && y_pointer == 28)
||(x_pointer == 141 && y_pointer == 28)
||(x_pointer == 142 && y_pointer == 28)
||(x_pointer == 23 && y_pointer == 29)
||(x_pointer == 24 && y_pointer == 29)
||(x_pointer == 25 && y_pointer == 29)
||(x_pointer == 26 && y_pointer == 29)
||(x_pointer == 27 && y_pointer == 29)
||(x_pointer == 28 && y_pointer == 29)
||(x_pointer == 29 && y_pointer == 29)
||(x_pointer == 30 && y_pointer == 29)
||(x_pointer == 31 && y_pointer == 29)
||(x_pointer == 134 && y_pointer == 29)
||(x_pointer == 135 && y_pointer == 29)
||(x_pointer == 136 && y_pointer == 29)
||(x_pointer == 137 && y_pointer == 29)
||(x_pointer == 138 && y_pointer == 29)
||(x_pointer == 139 && y_pointer == 29)
||(x_pointer == 140 && y_pointer == 29)
||(x_pointer == 141 && y_pointer == 29)
||(x_pointer == 142 && y_pointer == 29)
||(x_pointer == 23 && y_pointer == 30)
||(x_pointer == 24 && y_pointer == 30)
||(x_pointer == 25 && y_pointer == 30)
||(x_pointer == 26 && y_pointer == 30)
||(x_pointer == 27 && y_pointer == 30)
||(x_pointer == 28 && y_pointer == 30)
||(x_pointer == 29 && y_pointer == 30)
||(x_pointer == 30 && y_pointer == 30)
||(x_pointer == 31 && y_pointer == 30)
||(x_pointer == 134 && y_pointer == 30)
||(x_pointer == 135 && y_pointer == 30)
||(x_pointer == 136 && y_pointer == 30)
||(x_pointer == 137 && y_pointer == 30)
||(x_pointer == 138 && y_pointer == 30)
||(x_pointer == 139 && y_pointer == 30)
||(x_pointer == 140 && y_pointer == 30)
||(x_pointer == 141 && y_pointer == 30)
||(x_pointer == 142 && y_pointer == 30)
||(x_pointer == 23 && y_pointer == 31)
||(x_pointer == 24 && y_pointer == 31)
||(x_pointer == 25 && y_pointer == 31)
||(x_pointer == 26 && y_pointer == 31)
||(x_pointer == 27 && y_pointer == 31)
||(x_pointer == 28 && y_pointer == 31)
||(x_pointer == 29 && y_pointer == 31)
||(x_pointer == 30 && y_pointer == 31)
||(x_pointer == 31 && y_pointer == 31)
||(x_pointer == 134 && y_pointer == 31)
||(x_pointer == 135 && y_pointer == 31)
||(x_pointer == 136 && y_pointer == 31)
||(x_pointer == 137 && y_pointer == 31)
||(x_pointer == 138 && y_pointer == 31)
||(x_pointer == 139 && y_pointer == 31)
||(x_pointer == 140 && y_pointer == 31)
||(x_pointer == 141 && y_pointer == 31)
||(x_pointer == 142 && y_pointer == 31)
||(x_pointer == 23 && y_pointer == 32)
||(x_pointer == 24 && y_pointer == 32)
||(x_pointer == 25 && y_pointer == 32)
||(x_pointer == 26 && y_pointer == 32)
||(x_pointer == 27 && y_pointer == 32)
||(x_pointer == 28 && y_pointer == 32)
||(x_pointer == 29 && y_pointer == 32)
||(x_pointer == 30 && y_pointer == 32)
||(x_pointer == 31 && y_pointer == 32)
||(x_pointer == 50 && y_pointer == 32)
||(x_pointer == 51 && y_pointer == 32)
||(x_pointer == 52 && y_pointer == 32)
||(x_pointer == 53 && y_pointer == 32)
||(x_pointer == 54 && y_pointer == 32)
||(x_pointer == 55 && y_pointer == 32)
||(x_pointer == 56 && y_pointer == 32)
||(x_pointer == 57 && y_pointer == 32)
||(x_pointer == 58 && y_pointer == 32)
||(x_pointer == 59 && y_pointer == 32)
||(x_pointer == 60 && y_pointer == 32)
||(x_pointer == 61 && y_pointer == 32)
||(x_pointer == 62 && y_pointer == 32)
||(x_pointer == 63 && y_pointer == 32)
||(x_pointer == 64 && y_pointer == 32)
||(x_pointer == 65 && y_pointer == 32)
||(x_pointer == 66 && y_pointer == 32)
||(x_pointer == 67 && y_pointer == 32)
||(x_pointer == 68 && y_pointer == 32)
||(x_pointer == 69 && y_pointer == 32)
||(x_pointer == 70 && y_pointer == 32)
||(x_pointer == 71 && y_pointer == 32)
||(x_pointer == 72 && y_pointer == 32)
||(x_pointer == 73 && y_pointer == 32)
||(x_pointer == 74 && y_pointer == 32)
||(x_pointer == 75 && y_pointer == 32)
||(x_pointer == 76 && y_pointer == 32)
||(x_pointer == 77 && y_pointer == 32)
||(x_pointer == 78 && y_pointer == 32)
||(x_pointer == 79 && y_pointer == 32)
||(x_pointer == 80 && y_pointer == 32)
||(x_pointer == 81 && y_pointer == 32)
||(x_pointer == 82 && y_pointer == 32)
||(x_pointer == 83 && y_pointer == 32)
||(x_pointer == 84 && y_pointer == 32)
||(x_pointer == 85 && y_pointer == 32)
||(x_pointer == 86 && y_pointer == 32)
||(x_pointer == 87 && y_pointer == 32)
||(x_pointer == 88 && y_pointer == 32)
||(x_pointer == 89 && y_pointer == 32)
||(x_pointer == 90 && y_pointer == 32)
||(x_pointer == 91 && y_pointer == 32)
||(x_pointer == 92 && y_pointer == 32)
||(x_pointer == 93 && y_pointer == 32)
||(x_pointer == 94 && y_pointer == 32)
||(x_pointer == 95 && y_pointer == 32)
||(x_pointer == 96 && y_pointer == 32)
||(x_pointer == 97 && y_pointer == 32)
||(x_pointer == 98 && y_pointer == 32)
||(x_pointer == 99 && y_pointer == 32)
||(x_pointer == 100 && y_pointer == 32)
||(x_pointer == 101 && y_pointer == 32)
||(x_pointer == 102 && y_pointer == 32)
||(x_pointer == 103 && y_pointer == 32)
||(x_pointer == 104 && y_pointer == 32)
||(x_pointer == 105 && y_pointer == 32)
||(x_pointer == 106 && y_pointer == 32)
||(x_pointer == 107 && y_pointer == 32)
||(x_pointer == 108 && y_pointer == 32)
||(x_pointer == 109 && y_pointer == 32)
||(x_pointer == 110 && y_pointer == 32)
||(x_pointer == 111 && y_pointer == 32)
||(x_pointer == 112 && y_pointer == 32)
||(x_pointer == 113 && y_pointer == 32)
||(x_pointer == 114 && y_pointer == 32)
||(x_pointer == 115 && y_pointer == 32)
||(x_pointer == 134 && y_pointer == 32)
||(x_pointer == 135 && y_pointer == 32)
||(x_pointer == 136 && y_pointer == 32)
||(x_pointer == 137 && y_pointer == 32)
||(x_pointer == 138 && y_pointer == 32)
||(x_pointer == 139 && y_pointer == 32)
||(x_pointer == 140 && y_pointer == 32)
||(x_pointer == 141 && y_pointer == 32)
||(x_pointer == 142 && y_pointer == 32)
||(x_pointer == 23 && y_pointer == 33)
||(x_pointer == 24 && y_pointer == 33)
||(x_pointer == 25 && y_pointer == 33)
||(x_pointer == 26 && y_pointer == 33)
||(x_pointer == 27 && y_pointer == 33)
||(x_pointer == 28 && y_pointer == 33)
||(x_pointer == 29 && y_pointer == 33)
||(x_pointer == 30 && y_pointer == 33)
||(x_pointer == 31 && y_pointer == 33)
||(x_pointer == 50 && y_pointer == 33)
||(x_pointer == 51 && y_pointer == 33)
||(x_pointer == 52 && y_pointer == 33)
||(x_pointer == 53 && y_pointer == 33)
||(x_pointer == 54 && y_pointer == 33)
||(x_pointer == 55 && y_pointer == 33)
||(x_pointer == 56 && y_pointer == 33)
||(x_pointer == 57 && y_pointer == 33)
||(x_pointer == 58 && y_pointer == 33)
||(x_pointer == 59 && y_pointer == 33)
||(x_pointer == 60 && y_pointer == 33)
||(x_pointer == 61 && y_pointer == 33)
||(x_pointer == 62 && y_pointer == 33)
||(x_pointer == 63 && y_pointer == 33)
||(x_pointer == 64 && y_pointer == 33)
||(x_pointer == 65 && y_pointer == 33)
||(x_pointer == 66 && y_pointer == 33)
||(x_pointer == 67 && y_pointer == 33)
||(x_pointer == 68 && y_pointer == 33)
||(x_pointer == 69 && y_pointer == 33)
||(x_pointer == 70 && y_pointer == 33)
||(x_pointer == 71 && y_pointer == 33)
||(x_pointer == 72 && y_pointer == 33)
||(x_pointer == 73 && y_pointer == 33)
||(x_pointer == 74 && y_pointer == 33)
||(x_pointer == 75 && y_pointer == 33)
||(x_pointer == 76 && y_pointer == 33)
||(x_pointer == 77 && y_pointer == 33)
||(x_pointer == 78 && y_pointer == 33)
||(x_pointer == 79 && y_pointer == 33)
||(x_pointer == 80 && y_pointer == 33)
||(x_pointer == 81 && y_pointer == 33)
||(x_pointer == 82 && y_pointer == 33)
||(x_pointer == 83 && y_pointer == 33)
||(x_pointer == 84 && y_pointer == 33)
||(x_pointer == 85 && y_pointer == 33)
||(x_pointer == 86 && y_pointer == 33)
||(x_pointer == 87 && y_pointer == 33)
||(x_pointer == 88 && y_pointer == 33)
||(x_pointer == 89 && y_pointer == 33)
||(x_pointer == 90 && y_pointer == 33)
||(x_pointer == 91 && y_pointer == 33)
||(x_pointer == 92 && y_pointer == 33)
||(x_pointer == 93 && y_pointer == 33)
||(x_pointer == 94 && y_pointer == 33)
||(x_pointer == 95 && y_pointer == 33)
||(x_pointer == 96 && y_pointer == 33)
||(x_pointer == 97 && y_pointer == 33)
||(x_pointer == 98 && y_pointer == 33)
||(x_pointer == 99 && y_pointer == 33)
||(x_pointer == 100 && y_pointer == 33)
||(x_pointer == 101 && y_pointer == 33)
||(x_pointer == 102 && y_pointer == 33)
||(x_pointer == 103 && y_pointer == 33)
||(x_pointer == 104 && y_pointer == 33)
||(x_pointer == 105 && y_pointer == 33)
||(x_pointer == 106 && y_pointer == 33)
||(x_pointer == 107 && y_pointer == 33)
||(x_pointer == 108 && y_pointer == 33)
||(x_pointer == 109 && y_pointer == 33)
||(x_pointer == 110 && y_pointer == 33)
||(x_pointer == 111 && y_pointer == 33)
||(x_pointer == 112 && y_pointer == 33)
||(x_pointer == 113 && y_pointer == 33)
||(x_pointer == 114 && y_pointer == 33)
||(x_pointer == 115 && y_pointer == 33)
||(x_pointer == 134 && y_pointer == 33)
||(x_pointer == 135 && y_pointer == 33)
||(x_pointer == 136 && y_pointer == 33)
||(x_pointer == 137 && y_pointer == 33)
||(x_pointer == 138 && y_pointer == 33)
||(x_pointer == 139 && y_pointer == 33)
||(x_pointer == 140 && y_pointer == 33)
||(x_pointer == 141 && y_pointer == 33)
||(x_pointer == 142 && y_pointer == 33)
||(x_pointer == 23 && y_pointer == 34)
||(x_pointer == 24 && y_pointer == 34)
||(x_pointer == 25 && y_pointer == 34)
||(x_pointer == 26 && y_pointer == 34)
||(x_pointer == 27 && y_pointer == 34)
||(x_pointer == 28 && y_pointer == 34)
||(x_pointer == 29 && y_pointer == 34)
||(x_pointer == 30 && y_pointer == 34)
||(x_pointer == 31 && y_pointer == 34)
||(x_pointer == 50 && y_pointer == 34)
||(x_pointer == 51 && y_pointer == 34)
||(x_pointer == 52 && y_pointer == 34)
||(x_pointer == 53 && y_pointer == 34)
||(x_pointer == 54 && y_pointer == 34)
||(x_pointer == 55 && y_pointer == 34)
||(x_pointer == 56 && y_pointer == 34)
||(x_pointer == 57 && y_pointer == 34)
||(x_pointer == 58 && y_pointer == 34)
||(x_pointer == 59 && y_pointer == 34)
||(x_pointer == 60 && y_pointer == 34)
||(x_pointer == 61 && y_pointer == 34)
||(x_pointer == 62 && y_pointer == 34)
||(x_pointer == 63 && y_pointer == 34)
||(x_pointer == 64 && y_pointer == 34)
||(x_pointer == 65 && y_pointer == 34)
||(x_pointer == 66 && y_pointer == 34)
||(x_pointer == 67 && y_pointer == 34)
||(x_pointer == 68 && y_pointer == 34)
||(x_pointer == 69 && y_pointer == 34)
||(x_pointer == 70 && y_pointer == 34)
||(x_pointer == 71 && y_pointer == 34)
||(x_pointer == 72 && y_pointer == 34)
||(x_pointer == 73 && y_pointer == 34)
||(x_pointer == 74 && y_pointer == 34)
||(x_pointer == 75 && y_pointer == 34)
||(x_pointer == 76 && y_pointer == 34)
||(x_pointer == 77 && y_pointer == 34)
||(x_pointer == 78 && y_pointer == 34)
||(x_pointer == 79 && y_pointer == 34)
||(x_pointer == 80 && y_pointer == 34)
||(x_pointer == 81 && y_pointer == 34)
||(x_pointer == 82 && y_pointer == 34)
||(x_pointer == 83 && y_pointer == 34)
||(x_pointer == 84 && y_pointer == 34)
||(x_pointer == 85 && y_pointer == 34)
||(x_pointer == 86 && y_pointer == 34)
||(x_pointer == 87 && y_pointer == 34)
||(x_pointer == 88 && y_pointer == 34)
||(x_pointer == 89 && y_pointer == 34)
||(x_pointer == 90 && y_pointer == 34)
||(x_pointer == 91 && y_pointer == 34)
||(x_pointer == 92 && y_pointer == 34)
||(x_pointer == 93 && y_pointer == 34)
||(x_pointer == 94 && y_pointer == 34)
||(x_pointer == 95 && y_pointer == 34)
||(x_pointer == 96 && y_pointer == 34)
||(x_pointer == 97 && y_pointer == 34)
||(x_pointer == 98 && y_pointer == 34)
||(x_pointer == 99 && y_pointer == 34)
||(x_pointer == 100 && y_pointer == 34)
||(x_pointer == 101 && y_pointer == 34)
||(x_pointer == 102 && y_pointer == 34)
||(x_pointer == 103 && y_pointer == 34)
||(x_pointer == 104 && y_pointer == 34)
||(x_pointer == 105 && y_pointer == 34)
||(x_pointer == 106 && y_pointer == 34)
||(x_pointer == 107 && y_pointer == 34)
||(x_pointer == 108 && y_pointer == 34)
||(x_pointer == 109 && y_pointer == 34)
||(x_pointer == 110 && y_pointer == 34)
||(x_pointer == 111 && y_pointer == 34)
||(x_pointer == 112 && y_pointer == 34)
||(x_pointer == 113 && y_pointer == 34)
||(x_pointer == 114 && y_pointer == 34)
||(x_pointer == 115 && y_pointer == 34)
||(x_pointer == 134 && y_pointer == 34)
||(x_pointer == 135 && y_pointer == 34)
||(x_pointer == 136 && y_pointer == 34)
||(x_pointer == 137 && y_pointer == 34)
||(x_pointer == 138 && y_pointer == 34)
||(x_pointer == 139 && y_pointer == 34)
||(x_pointer == 140 && y_pointer == 34)
||(x_pointer == 141 && y_pointer == 34)
||(x_pointer == 142 && y_pointer == 34)
||(x_pointer == 23 && y_pointer == 35)
||(x_pointer == 24 && y_pointer == 35)
||(x_pointer == 25 && y_pointer == 35)
||(x_pointer == 26 && y_pointer == 35)
||(x_pointer == 27 && y_pointer == 35)
||(x_pointer == 28 && y_pointer == 35)
||(x_pointer == 29 && y_pointer == 35)
||(x_pointer == 30 && y_pointer == 35)
||(x_pointer == 31 && y_pointer == 35)
||(x_pointer == 50 && y_pointer == 35)
||(x_pointer == 51 && y_pointer == 35)
||(x_pointer == 52 && y_pointer == 35)
||(x_pointer == 53 && y_pointer == 35)
||(x_pointer == 54 && y_pointer == 35)
||(x_pointer == 55 && y_pointer == 35)
||(x_pointer == 56 && y_pointer == 35)
||(x_pointer == 57 && y_pointer == 35)
||(x_pointer == 58 && y_pointer == 35)
||(x_pointer == 59 && y_pointer == 35)
||(x_pointer == 60 && y_pointer == 35)
||(x_pointer == 61 && y_pointer == 35)
||(x_pointer == 62 && y_pointer == 35)
||(x_pointer == 63 && y_pointer == 35)
||(x_pointer == 64 && y_pointer == 35)
||(x_pointer == 65 && y_pointer == 35)
||(x_pointer == 66 && y_pointer == 35)
||(x_pointer == 67 && y_pointer == 35)
||(x_pointer == 68 && y_pointer == 35)
||(x_pointer == 69 && y_pointer == 35)
||(x_pointer == 70 && y_pointer == 35)
||(x_pointer == 71 && y_pointer == 35)
||(x_pointer == 72 && y_pointer == 35)
||(x_pointer == 73 && y_pointer == 35)
||(x_pointer == 74 && y_pointer == 35)
||(x_pointer == 75 && y_pointer == 35)
||(x_pointer == 76 && y_pointer == 35)
||(x_pointer == 77 && y_pointer == 35)
||(x_pointer == 78 && y_pointer == 35)
||(x_pointer == 79 && y_pointer == 35)
||(x_pointer == 80 && y_pointer == 35)
||(x_pointer == 81 && y_pointer == 35)
||(x_pointer == 82 && y_pointer == 35)
||(x_pointer == 83 && y_pointer == 35)
||(x_pointer == 84 && y_pointer == 35)
||(x_pointer == 85 && y_pointer == 35)
||(x_pointer == 86 && y_pointer == 35)
||(x_pointer == 87 && y_pointer == 35)
||(x_pointer == 88 && y_pointer == 35)
||(x_pointer == 89 && y_pointer == 35)
||(x_pointer == 90 && y_pointer == 35)
||(x_pointer == 91 && y_pointer == 35)
||(x_pointer == 92 && y_pointer == 35)
||(x_pointer == 93 && y_pointer == 35)
||(x_pointer == 94 && y_pointer == 35)
||(x_pointer == 95 && y_pointer == 35)
||(x_pointer == 96 && y_pointer == 35)
||(x_pointer == 97 && y_pointer == 35)
||(x_pointer == 98 && y_pointer == 35)
||(x_pointer == 99 && y_pointer == 35)
||(x_pointer == 100 && y_pointer == 35)
||(x_pointer == 101 && y_pointer == 35)
||(x_pointer == 102 && y_pointer == 35)
||(x_pointer == 103 && y_pointer == 35)
||(x_pointer == 104 && y_pointer == 35)
||(x_pointer == 105 && y_pointer == 35)
||(x_pointer == 106 && y_pointer == 35)
||(x_pointer == 107 && y_pointer == 35)
||(x_pointer == 108 && y_pointer == 35)
||(x_pointer == 109 && y_pointer == 35)
||(x_pointer == 110 && y_pointer == 35)
||(x_pointer == 111 && y_pointer == 35)
||(x_pointer == 112 && y_pointer == 35)
||(x_pointer == 113 && y_pointer == 35)
||(x_pointer == 114 && y_pointer == 35)
||(x_pointer == 115 && y_pointer == 35)
||(x_pointer == 134 && y_pointer == 35)
||(x_pointer == 135 && y_pointer == 35)
||(x_pointer == 136 && y_pointer == 35)
||(x_pointer == 137 && y_pointer == 35)
||(x_pointer == 138 && y_pointer == 35)
||(x_pointer == 139 && y_pointer == 35)
||(x_pointer == 140 && y_pointer == 35)
||(x_pointer == 141 && y_pointer == 35)
||(x_pointer == 142 && y_pointer == 35)
||(x_pointer == 23 && y_pointer == 36)
||(x_pointer == 24 && y_pointer == 36)
||(x_pointer == 25 && y_pointer == 36)
||(x_pointer == 26 && y_pointer == 36)
||(x_pointer == 27 && y_pointer == 36)
||(x_pointer == 28 && y_pointer == 36)
||(x_pointer == 29 && y_pointer == 36)
||(x_pointer == 30 && y_pointer == 36)
||(x_pointer == 31 && y_pointer == 36)
||(x_pointer == 50 && y_pointer == 36)
||(x_pointer == 51 && y_pointer == 36)
||(x_pointer == 52 && y_pointer == 36)
||(x_pointer == 53 && y_pointer == 36)
||(x_pointer == 54 && y_pointer == 36)
||(x_pointer == 55 && y_pointer == 36)
||(x_pointer == 56 && y_pointer == 36)
||(x_pointer == 57 && y_pointer == 36)
||(x_pointer == 58 && y_pointer == 36)
||(x_pointer == 59 && y_pointer == 36)
||(x_pointer == 60 && y_pointer == 36)
||(x_pointer == 61 && y_pointer == 36)
||(x_pointer == 62 && y_pointer == 36)
||(x_pointer == 63 && y_pointer == 36)
||(x_pointer == 64 && y_pointer == 36)
||(x_pointer == 65 && y_pointer == 36)
||(x_pointer == 66 && y_pointer == 36)
||(x_pointer == 67 && y_pointer == 36)
||(x_pointer == 68 && y_pointer == 36)
||(x_pointer == 69 && y_pointer == 36)
||(x_pointer == 70 && y_pointer == 36)
||(x_pointer == 71 && y_pointer == 36)
||(x_pointer == 72 && y_pointer == 36)
||(x_pointer == 73 && y_pointer == 36)
||(x_pointer == 74 && y_pointer == 36)
||(x_pointer == 75 && y_pointer == 36)
||(x_pointer == 76 && y_pointer == 36)
||(x_pointer == 77 && y_pointer == 36)
||(x_pointer == 78 && y_pointer == 36)
||(x_pointer == 79 && y_pointer == 36)
||(x_pointer == 80 && y_pointer == 36)
||(x_pointer == 81 && y_pointer == 36)
||(x_pointer == 82 && y_pointer == 36)
||(x_pointer == 83 && y_pointer == 36)
||(x_pointer == 84 && y_pointer == 36)
||(x_pointer == 85 && y_pointer == 36)
||(x_pointer == 86 && y_pointer == 36)
||(x_pointer == 87 && y_pointer == 36)
||(x_pointer == 88 && y_pointer == 36)
||(x_pointer == 89 && y_pointer == 36)
||(x_pointer == 90 && y_pointer == 36)
||(x_pointer == 91 && y_pointer == 36)
||(x_pointer == 92 && y_pointer == 36)
||(x_pointer == 93 && y_pointer == 36)
||(x_pointer == 94 && y_pointer == 36)
||(x_pointer == 95 && y_pointer == 36)
||(x_pointer == 96 && y_pointer == 36)
||(x_pointer == 97 && y_pointer == 36)
||(x_pointer == 98 && y_pointer == 36)
||(x_pointer == 99 && y_pointer == 36)
||(x_pointer == 100 && y_pointer == 36)
||(x_pointer == 101 && y_pointer == 36)
||(x_pointer == 102 && y_pointer == 36)
||(x_pointer == 103 && y_pointer == 36)
||(x_pointer == 104 && y_pointer == 36)
||(x_pointer == 105 && y_pointer == 36)
||(x_pointer == 106 && y_pointer == 36)
||(x_pointer == 107 && y_pointer == 36)
||(x_pointer == 108 && y_pointer == 36)
||(x_pointer == 109 && y_pointer == 36)
||(x_pointer == 110 && y_pointer == 36)
||(x_pointer == 111 && y_pointer == 36)
||(x_pointer == 112 && y_pointer == 36)
||(x_pointer == 113 && y_pointer == 36)
||(x_pointer == 114 && y_pointer == 36)
||(x_pointer == 115 && y_pointer == 36)
||(x_pointer == 134 && y_pointer == 36)
||(x_pointer == 135 && y_pointer == 36)
||(x_pointer == 136 && y_pointer == 36)
||(x_pointer == 137 && y_pointer == 36)
||(x_pointer == 138 && y_pointer == 36)
||(x_pointer == 139 && y_pointer == 36)
||(x_pointer == 140 && y_pointer == 36)
||(x_pointer == 141 && y_pointer == 36)
||(x_pointer == 142 && y_pointer == 36)
||(x_pointer == 50 && y_pointer == 37)
||(x_pointer == 51 && y_pointer == 37)
||(x_pointer == 52 && y_pointer == 37)
||(x_pointer == 53 && y_pointer == 37)
||(x_pointer == 54 && y_pointer == 37)
||(x_pointer == 55 && y_pointer == 37)
||(x_pointer == 56 && y_pointer == 37)
||(x_pointer == 57 && y_pointer == 37)
||(x_pointer == 58 && y_pointer == 37)
||(x_pointer == 59 && y_pointer == 37)
||(x_pointer == 60 && y_pointer == 37)
||(x_pointer == 61 && y_pointer == 37)
||(x_pointer == 62 && y_pointer == 37)
||(x_pointer == 63 && y_pointer == 37)
||(x_pointer == 64 && y_pointer == 37)
||(x_pointer == 65 && y_pointer == 37)
||(x_pointer == 66 && y_pointer == 37)
||(x_pointer == 67 && y_pointer == 37)
||(x_pointer == 68 && y_pointer == 37)
||(x_pointer == 69 && y_pointer == 37)
||(x_pointer == 70 && y_pointer == 37)
||(x_pointer == 71 && y_pointer == 37)
||(x_pointer == 72 && y_pointer == 37)
||(x_pointer == 73 && y_pointer == 37)
||(x_pointer == 74 && y_pointer == 37)
||(x_pointer == 75 && y_pointer == 37)
||(x_pointer == 76 && y_pointer == 37)
||(x_pointer == 77 && y_pointer == 37)
||(x_pointer == 78 && y_pointer == 37)
||(x_pointer == 79 && y_pointer == 37)
||(x_pointer == 80 && y_pointer == 37)
||(x_pointer == 81 && y_pointer == 37)
||(x_pointer == 82 && y_pointer == 37)
||(x_pointer == 83 && y_pointer == 37)
||(x_pointer == 84 && y_pointer == 37)
||(x_pointer == 85 && y_pointer == 37)
||(x_pointer == 86 && y_pointer == 37)
||(x_pointer == 87 && y_pointer == 37)
||(x_pointer == 88 && y_pointer == 37)
||(x_pointer == 89 && y_pointer == 37)
||(x_pointer == 90 && y_pointer == 37)
||(x_pointer == 91 && y_pointer == 37)
||(x_pointer == 92 && y_pointer == 37)
||(x_pointer == 93 && y_pointer == 37)
||(x_pointer == 94 && y_pointer == 37)
||(x_pointer == 95 && y_pointer == 37)
||(x_pointer == 96 && y_pointer == 37)
||(x_pointer == 97 && y_pointer == 37)
||(x_pointer == 98 && y_pointer == 37)
||(x_pointer == 99 && y_pointer == 37)
||(x_pointer == 100 && y_pointer == 37)
||(x_pointer == 101 && y_pointer == 37)
||(x_pointer == 102 && y_pointer == 37)
||(x_pointer == 103 && y_pointer == 37)
||(x_pointer == 104 && y_pointer == 37)
||(x_pointer == 105 && y_pointer == 37)
||(x_pointer == 106 && y_pointer == 37)
||(x_pointer == 107 && y_pointer == 37)
||(x_pointer == 108 && y_pointer == 37)
||(x_pointer == 109 && y_pointer == 37)
||(x_pointer == 110 && y_pointer == 37)
||(x_pointer == 111 && y_pointer == 37)
||(x_pointer == 112 && y_pointer == 37)
||(x_pointer == 113 && y_pointer == 37)
||(x_pointer == 114 && y_pointer == 37)
||(x_pointer == 115 && y_pointer == 37)
||(x_pointer == 50 && y_pointer == 38)
||(x_pointer == 51 && y_pointer == 38)
||(x_pointer == 52 && y_pointer == 38)
||(x_pointer == 53 && y_pointer == 38)
||(x_pointer == 54 && y_pointer == 38)
||(x_pointer == 55 && y_pointer == 38)
||(x_pointer == 56 && y_pointer == 38)
||(x_pointer == 57 && y_pointer == 38)
||(x_pointer == 58 && y_pointer == 38)
||(x_pointer == 59 && y_pointer == 38)
||(x_pointer == 60 && y_pointer == 38)
||(x_pointer == 61 && y_pointer == 38)
||(x_pointer == 62 && y_pointer == 38)
||(x_pointer == 63 && y_pointer == 38)
||(x_pointer == 64 && y_pointer == 38)
||(x_pointer == 65 && y_pointer == 38)
||(x_pointer == 66 && y_pointer == 38)
||(x_pointer == 67 && y_pointer == 38)
||(x_pointer == 68 && y_pointer == 38)
||(x_pointer == 69 && y_pointer == 38)
||(x_pointer == 70 && y_pointer == 38)
||(x_pointer == 71 && y_pointer == 38)
||(x_pointer == 72 && y_pointer == 38)
||(x_pointer == 73 && y_pointer == 38)
||(x_pointer == 74 && y_pointer == 38)
||(x_pointer == 75 && y_pointer == 38)
||(x_pointer == 76 && y_pointer == 38)
||(x_pointer == 77 && y_pointer == 38)
||(x_pointer == 78 && y_pointer == 38)
||(x_pointer == 79 && y_pointer == 38)
||(x_pointer == 80 && y_pointer == 38)
||(x_pointer == 81 && y_pointer == 38)
||(x_pointer == 82 && y_pointer == 38)
||(x_pointer == 83 && y_pointer == 38)
||(x_pointer == 84 && y_pointer == 38)
||(x_pointer == 85 && y_pointer == 38)
||(x_pointer == 86 && y_pointer == 38)
||(x_pointer == 87 && y_pointer == 38)
||(x_pointer == 88 && y_pointer == 38)
||(x_pointer == 89 && y_pointer == 38)
||(x_pointer == 90 && y_pointer == 38)
||(x_pointer == 91 && y_pointer == 38)
||(x_pointer == 92 && y_pointer == 38)
||(x_pointer == 93 && y_pointer == 38)
||(x_pointer == 94 && y_pointer == 38)
||(x_pointer == 95 && y_pointer == 38)
||(x_pointer == 96 && y_pointer == 38)
||(x_pointer == 97 && y_pointer == 38)
||(x_pointer == 98 && y_pointer == 38)
||(x_pointer == 99 && y_pointer == 38)
||(x_pointer == 100 && y_pointer == 38)
||(x_pointer == 101 && y_pointer == 38)
||(x_pointer == 102 && y_pointer == 38)
||(x_pointer == 103 && y_pointer == 38)
||(x_pointer == 104 && y_pointer == 38)
||(x_pointer == 105 && y_pointer == 38)
||(x_pointer == 106 && y_pointer == 38)
||(x_pointer == 107 && y_pointer == 38)
||(x_pointer == 108 && y_pointer == 38)
||(x_pointer == 109 && y_pointer == 38)
||(x_pointer == 110 && y_pointer == 38)
||(x_pointer == 111 && y_pointer == 38)
||(x_pointer == 112 && y_pointer == 38)
||(x_pointer == 113 && y_pointer == 38)
||(x_pointer == 114 && y_pointer == 38)
||(x_pointer == 115 && y_pointer == 38)
||(x_pointer == 50 && y_pointer == 39)
||(x_pointer == 51 && y_pointer == 39)
||(x_pointer == 52 && y_pointer == 39)
||(x_pointer == 53 && y_pointer == 39)
||(x_pointer == 54 && y_pointer == 39)
||(x_pointer == 55 && y_pointer == 39)
||(x_pointer == 56 && y_pointer == 39)
||(x_pointer == 57 && y_pointer == 39)
||(x_pointer == 58 && y_pointer == 39)
||(x_pointer == 59 && y_pointer == 39)
||(x_pointer == 60 && y_pointer == 39)
||(x_pointer == 61 && y_pointer == 39)
||(x_pointer == 62 && y_pointer == 39)
||(x_pointer == 63 && y_pointer == 39)
||(x_pointer == 64 && y_pointer == 39)
||(x_pointer == 65 && y_pointer == 39)
||(x_pointer == 66 && y_pointer == 39)
||(x_pointer == 67 && y_pointer == 39)
||(x_pointer == 68 && y_pointer == 39)
||(x_pointer == 69 && y_pointer == 39)
||(x_pointer == 70 && y_pointer == 39)
||(x_pointer == 71 && y_pointer == 39)
||(x_pointer == 72 && y_pointer == 39)
||(x_pointer == 73 && y_pointer == 39)
||(x_pointer == 74 && y_pointer == 39)
||(x_pointer == 75 && y_pointer == 39)
||(x_pointer == 76 && y_pointer == 39)
||(x_pointer == 77 && y_pointer == 39)
||(x_pointer == 78 && y_pointer == 39)
||(x_pointer == 79 && y_pointer == 39)
||(x_pointer == 80 && y_pointer == 39)
||(x_pointer == 81 && y_pointer == 39)
||(x_pointer == 82 && y_pointer == 39)
||(x_pointer == 83 && y_pointer == 39)
||(x_pointer == 84 && y_pointer == 39)
||(x_pointer == 85 && y_pointer == 39)
||(x_pointer == 86 && y_pointer == 39)
||(x_pointer == 87 && y_pointer == 39)
||(x_pointer == 88 && y_pointer == 39)
||(x_pointer == 89 && y_pointer == 39)
||(x_pointer == 90 && y_pointer == 39)
||(x_pointer == 91 && y_pointer == 39)
||(x_pointer == 92 && y_pointer == 39)
||(x_pointer == 93 && y_pointer == 39)
||(x_pointer == 94 && y_pointer == 39)
||(x_pointer == 95 && y_pointer == 39)
||(x_pointer == 96 && y_pointer == 39)
||(x_pointer == 97 && y_pointer == 39)
||(x_pointer == 98 && y_pointer == 39)
||(x_pointer == 99 && y_pointer == 39)
||(x_pointer == 100 && y_pointer == 39)
||(x_pointer == 101 && y_pointer == 39)
||(x_pointer == 102 && y_pointer == 39)
||(x_pointer == 103 && y_pointer == 39)
||(x_pointer == 104 && y_pointer == 39)
||(x_pointer == 105 && y_pointer == 39)
||(x_pointer == 106 && y_pointer == 39)
||(x_pointer == 107 && y_pointer == 39)
||(x_pointer == 108 && y_pointer == 39)
||(x_pointer == 109 && y_pointer == 39)
||(x_pointer == 110 && y_pointer == 39)
||(x_pointer == 111 && y_pointer == 39)
||(x_pointer == 112 && y_pointer == 39)
||(x_pointer == 113 && y_pointer == 39)
||(x_pointer == 114 && y_pointer == 39)
||(x_pointer == 115 && y_pointer == 39)
||(x_pointer == 50 && y_pointer == 40)
||(x_pointer == 51 && y_pointer == 40)
||(x_pointer == 52 && y_pointer == 40)
||(x_pointer == 53 && y_pointer == 40)
||(x_pointer == 54 && y_pointer == 40)
||(x_pointer == 55 && y_pointer == 40)
||(x_pointer == 56 && y_pointer == 40)
||(x_pointer == 57 && y_pointer == 40)
||(x_pointer == 58 && y_pointer == 40)
||(x_pointer == 59 && y_pointer == 40)
||(x_pointer == 60 && y_pointer == 40)
||(x_pointer == 61 && y_pointer == 40)
||(x_pointer == 62 && y_pointer == 40)
||(x_pointer == 63 && y_pointer == 40)
||(x_pointer == 64 && y_pointer == 40)
||(x_pointer == 65 && y_pointer == 40)
||(x_pointer == 66 && y_pointer == 40)
||(x_pointer == 67 && y_pointer == 40)
||(x_pointer == 68 && y_pointer == 40)
||(x_pointer == 69 && y_pointer == 40)
||(x_pointer == 70 && y_pointer == 40)
||(x_pointer == 71 && y_pointer == 40)
||(x_pointer == 72 && y_pointer == 40)
||(x_pointer == 73 && y_pointer == 40)
||(x_pointer == 74 && y_pointer == 40)
||(x_pointer == 75 && y_pointer == 40)
||(x_pointer == 76 && y_pointer == 40)
||(x_pointer == 77 && y_pointer == 40)
||(x_pointer == 78 && y_pointer == 40)
||(x_pointer == 79 && y_pointer == 40)
||(x_pointer == 80 && y_pointer == 40)
||(x_pointer == 81 && y_pointer == 40)
||(x_pointer == 82 && y_pointer == 40)
||(x_pointer == 83 && y_pointer == 40)
||(x_pointer == 84 && y_pointer == 40)
||(x_pointer == 85 && y_pointer == 40)
||(x_pointer == 86 && y_pointer == 40)
||(x_pointer == 87 && y_pointer == 40)
||(x_pointer == 88 && y_pointer == 40)
||(x_pointer == 89 && y_pointer == 40)
||(x_pointer == 90 && y_pointer == 40)
||(x_pointer == 91 && y_pointer == 40)
||(x_pointer == 92 && y_pointer == 40)
||(x_pointer == 93 && y_pointer == 40)
||(x_pointer == 94 && y_pointer == 40)
||(x_pointer == 95 && y_pointer == 40)
||(x_pointer == 96 && y_pointer == 40)
||(x_pointer == 97 && y_pointer == 40)
||(x_pointer == 98 && y_pointer == 40)
||(x_pointer == 99 && y_pointer == 40)
||(x_pointer == 100 && y_pointer == 40)
||(x_pointer == 101 && y_pointer == 40)
||(x_pointer == 102 && y_pointer == 40)
||(x_pointer == 103 && y_pointer == 40)
||(x_pointer == 104 && y_pointer == 40)
||(x_pointer == 105 && y_pointer == 40)
||(x_pointer == 106 && y_pointer == 40)
||(x_pointer == 107 && y_pointer == 40)
||(x_pointer == 108 && y_pointer == 40)
||(x_pointer == 109 && y_pointer == 40)
||(x_pointer == 110 && y_pointer == 40)
||(x_pointer == 111 && y_pointer == 40)
||(x_pointer == 112 && y_pointer == 40)
||(x_pointer == 113 && y_pointer == 40)
||(x_pointer == 114 && y_pointer == 40)
||(x_pointer == 115 && y_pointer == 40)
||(x_pointer == 50 && y_pointer == 68)
||(x_pointer == 51 && y_pointer == 68)
||(x_pointer == 52 && y_pointer == 68)
||(x_pointer == 53 && y_pointer == 68)
||(x_pointer == 54 && y_pointer == 68)
||(x_pointer == 55 && y_pointer == 68)
||(x_pointer == 56 && y_pointer == 68)
||(x_pointer == 57 && y_pointer == 68)
||(x_pointer == 58 && y_pointer == 68)
||(x_pointer == 59 && y_pointer == 68)
||(x_pointer == 60 && y_pointer == 68)
||(x_pointer == 61 && y_pointer == 68)
||(x_pointer == 62 && y_pointer == 68)
||(x_pointer == 63 && y_pointer == 68)
||(x_pointer == 64 && y_pointer == 68)
||(x_pointer == 65 && y_pointer == 68)
||(x_pointer == 66 && y_pointer == 68)
||(x_pointer == 67 && y_pointer == 68)
||(x_pointer == 68 && y_pointer == 68)
||(x_pointer == 69 && y_pointer == 68)
||(x_pointer == 70 && y_pointer == 68)
||(x_pointer == 71 && y_pointer == 68)
||(x_pointer == 72 && y_pointer == 68)
||(x_pointer == 73 && y_pointer == 68)
||(x_pointer == 74 && y_pointer == 68)
||(x_pointer == 75 && y_pointer == 68)
||(x_pointer == 76 && y_pointer == 68)
||(x_pointer == 77 && y_pointer == 68)
||(x_pointer == 78 && y_pointer == 68)
||(x_pointer == 79 && y_pointer == 68)
||(x_pointer == 80 && y_pointer == 68)
||(x_pointer == 81 && y_pointer == 68)
||(x_pointer == 82 && y_pointer == 68)
||(x_pointer == 83 && y_pointer == 68)
||(x_pointer == 84 && y_pointer == 68)
||(x_pointer == 85 && y_pointer == 68)
||(x_pointer == 86 && y_pointer == 68)
||(x_pointer == 87 && y_pointer == 68)
||(x_pointer == 88 && y_pointer == 68)
||(x_pointer == 89 && y_pointer == 68)
||(x_pointer == 90 && y_pointer == 68)
||(x_pointer == 91 && y_pointer == 68)
||(x_pointer == 92 && y_pointer == 68)
||(x_pointer == 93 && y_pointer == 68)
||(x_pointer == 94 && y_pointer == 68)
||(x_pointer == 95 && y_pointer == 68)
||(x_pointer == 96 && y_pointer == 68)
||(x_pointer == 97 && y_pointer == 68)
||(x_pointer == 98 && y_pointer == 68)
||(x_pointer == 99 && y_pointer == 68)
||(x_pointer == 100 && y_pointer == 68)
||(x_pointer == 101 && y_pointer == 68)
||(x_pointer == 102 && y_pointer == 68)
||(x_pointer == 103 && y_pointer == 68)
||(x_pointer == 104 && y_pointer == 68)
||(x_pointer == 105 && y_pointer == 68)
||(x_pointer == 106 && y_pointer == 68)
||(x_pointer == 107 && y_pointer == 68)
||(x_pointer == 108 && y_pointer == 68)
||(x_pointer == 109 && y_pointer == 68)
||(x_pointer == 110 && y_pointer == 68)
||(x_pointer == 111 && y_pointer == 68)
||(x_pointer == 112 && y_pointer == 68)
||(x_pointer == 113 && y_pointer == 68)
||(x_pointer == 114 && y_pointer == 68)
||(x_pointer == 115 && y_pointer == 68)
||(x_pointer == 50 && y_pointer == 69)
||(x_pointer == 51 && y_pointer == 69)
||(x_pointer == 52 && y_pointer == 69)
||(x_pointer == 53 && y_pointer == 69)
||(x_pointer == 54 && y_pointer == 69)
||(x_pointer == 55 && y_pointer == 69)
||(x_pointer == 56 && y_pointer == 69)
||(x_pointer == 57 && y_pointer == 69)
||(x_pointer == 58 && y_pointer == 69)
||(x_pointer == 59 && y_pointer == 69)
||(x_pointer == 60 && y_pointer == 69)
||(x_pointer == 61 && y_pointer == 69)
||(x_pointer == 62 && y_pointer == 69)
||(x_pointer == 63 && y_pointer == 69)
||(x_pointer == 64 && y_pointer == 69)
||(x_pointer == 65 && y_pointer == 69)
||(x_pointer == 66 && y_pointer == 69)
||(x_pointer == 67 && y_pointer == 69)
||(x_pointer == 68 && y_pointer == 69)
||(x_pointer == 69 && y_pointer == 69)
||(x_pointer == 70 && y_pointer == 69)
||(x_pointer == 71 && y_pointer == 69)
||(x_pointer == 72 && y_pointer == 69)
||(x_pointer == 73 && y_pointer == 69)
||(x_pointer == 74 && y_pointer == 69)
||(x_pointer == 75 && y_pointer == 69)
||(x_pointer == 76 && y_pointer == 69)
||(x_pointer == 77 && y_pointer == 69)
||(x_pointer == 78 && y_pointer == 69)
||(x_pointer == 79 && y_pointer == 69)
||(x_pointer == 80 && y_pointer == 69)
||(x_pointer == 81 && y_pointer == 69)
||(x_pointer == 82 && y_pointer == 69)
||(x_pointer == 83 && y_pointer == 69)
||(x_pointer == 84 && y_pointer == 69)
||(x_pointer == 85 && y_pointer == 69)
||(x_pointer == 86 && y_pointer == 69)
||(x_pointer == 87 && y_pointer == 69)
||(x_pointer == 88 && y_pointer == 69)
||(x_pointer == 89 && y_pointer == 69)
||(x_pointer == 90 && y_pointer == 69)
||(x_pointer == 91 && y_pointer == 69)
||(x_pointer == 92 && y_pointer == 69)
||(x_pointer == 93 && y_pointer == 69)
||(x_pointer == 94 && y_pointer == 69)
||(x_pointer == 95 && y_pointer == 69)
||(x_pointer == 96 && y_pointer == 69)
||(x_pointer == 97 && y_pointer == 69)
||(x_pointer == 98 && y_pointer == 69)
||(x_pointer == 99 && y_pointer == 69)
||(x_pointer == 100 && y_pointer == 69)
||(x_pointer == 101 && y_pointer == 69)
||(x_pointer == 102 && y_pointer == 69)
||(x_pointer == 103 && y_pointer == 69)
||(x_pointer == 104 && y_pointer == 69)
||(x_pointer == 105 && y_pointer == 69)
||(x_pointer == 106 && y_pointer == 69)
||(x_pointer == 107 && y_pointer == 69)
||(x_pointer == 108 && y_pointer == 69)
||(x_pointer == 109 && y_pointer == 69)
||(x_pointer == 110 && y_pointer == 69)
||(x_pointer == 111 && y_pointer == 69)
||(x_pointer == 112 && y_pointer == 69)
||(x_pointer == 113 && y_pointer == 69)
||(x_pointer == 114 && y_pointer == 69)
||(x_pointer == 115 && y_pointer == 69)
||(x_pointer == 50 && y_pointer == 70)
||(x_pointer == 51 && y_pointer == 70)
||(x_pointer == 52 && y_pointer == 70)
||(x_pointer == 53 && y_pointer == 70)
||(x_pointer == 54 && y_pointer == 70)
||(x_pointer == 55 && y_pointer == 70)
||(x_pointer == 56 && y_pointer == 70)
||(x_pointer == 57 && y_pointer == 70)
||(x_pointer == 58 && y_pointer == 70)
||(x_pointer == 59 && y_pointer == 70)
||(x_pointer == 60 && y_pointer == 70)
||(x_pointer == 61 && y_pointer == 70)
||(x_pointer == 62 && y_pointer == 70)
||(x_pointer == 63 && y_pointer == 70)
||(x_pointer == 64 && y_pointer == 70)
||(x_pointer == 65 && y_pointer == 70)
||(x_pointer == 66 && y_pointer == 70)
||(x_pointer == 67 && y_pointer == 70)
||(x_pointer == 68 && y_pointer == 70)
||(x_pointer == 69 && y_pointer == 70)
||(x_pointer == 70 && y_pointer == 70)
||(x_pointer == 71 && y_pointer == 70)
||(x_pointer == 72 && y_pointer == 70)
||(x_pointer == 73 && y_pointer == 70)
||(x_pointer == 74 && y_pointer == 70)
||(x_pointer == 75 && y_pointer == 70)
||(x_pointer == 76 && y_pointer == 70)
||(x_pointer == 77 && y_pointer == 70)
||(x_pointer == 78 && y_pointer == 70)
||(x_pointer == 79 && y_pointer == 70)
||(x_pointer == 80 && y_pointer == 70)
||(x_pointer == 81 && y_pointer == 70)
||(x_pointer == 82 && y_pointer == 70)
||(x_pointer == 83 && y_pointer == 70)
||(x_pointer == 84 && y_pointer == 70)
||(x_pointer == 85 && y_pointer == 70)
||(x_pointer == 86 && y_pointer == 70)
||(x_pointer == 87 && y_pointer == 70)
||(x_pointer == 88 && y_pointer == 70)
||(x_pointer == 89 && y_pointer == 70)
||(x_pointer == 90 && y_pointer == 70)
||(x_pointer == 91 && y_pointer == 70)
||(x_pointer == 92 && y_pointer == 70)
||(x_pointer == 93 && y_pointer == 70)
||(x_pointer == 94 && y_pointer == 70)
||(x_pointer == 95 && y_pointer == 70)
||(x_pointer == 96 && y_pointer == 70)
||(x_pointer == 97 && y_pointer == 70)
||(x_pointer == 98 && y_pointer == 70)
||(x_pointer == 99 && y_pointer == 70)
||(x_pointer == 100 && y_pointer == 70)
||(x_pointer == 101 && y_pointer == 70)
||(x_pointer == 102 && y_pointer == 70)
||(x_pointer == 103 && y_pointer == 70)
||(x_pointer == 104 && y_pointer == 70)
||(x_pointer == 105 && y_pointer == 70)
||(x_pointer == 106 && y_pointer == 70)
||(x_pointer == 107 && y_pointer == 70)
||(x_pointer == 108 && y_pointer == 70)
||(x_pointer == 109 && y_pointer == 70)
||(x_pointer == 110 && y_pointer == 70)
||(x_pointer == 111 && y_pointer == 70)
||(x_pointer == 112 && y_pointer == 70)
||(x_pointer == 113 && y_pointer == 70)
||(x_pointer == 114 && y_pointer == 70)
||(x_pointer == 115 && y_pointer == 70)
||(x_pointer == 50 && y_pointer == 71)
||(x_pointer == 51 && y_pointer == 71)
||(x_pointer == 52 && y_pointer == 71)
||(x_pointer == 53 && y_pointer == 71)
||(x_pointer == 54 && y_pointer == 71)
||(x_pointer == 55 && y_pointer == 71)
||(x_pointer == 56 && y_pointer == 71)
||(x_pointer == 57 && y_pointer == 71)
||(x_pointer == 58 && y_pointer == 71)
||(x_pointer == 59 && y_pointer == 71)
||(x_pointer == 60 && y_pointer == 71)
||(x_pointer == 61 && y_pointer == 71)
||(x_pointer == 62 && y_pointer == 71)
||(x_pointer == 63 && y_pointer == 71)
||(x_pointer == 64 && y_pointer == 71)
||(x_pointer == 65 && y_pointer == 71)
||(x_pointer == 66 && y_pointer == 71)
||(x_pointer == 67 && y_pointer == 71)
||(x_pointer == 68 && y_pointer == 71)
||(x_pointer == 69 && y_pointer == 71)
||(x_pointer == 70 && y_pointer == 71)
||(x_pointer == 71 && y_pointer == 71)
||(x_pointer == 72 && y_pointer == 71)
||(x_pointer == 73 && y_pointer == 71)
||(x_pointer == 74 && y_pointer == 71)
||(x_pointer == 75 && y_pointer == 71)
||(x_pointer == 76 && y_pointer == 71)
||(x_pointer == 77 && y_pointer == 71)
||(x_pointer == 78 && y_pointer == 71)
||(x_pointer == 79 && y_pointer == 71)
||(x_pointer == 80 && y_pointer == 71)
||(x_pointer == 81 && y_pointer == 71)
||(x_pointer == 82 && y_pointer == 71)
||(x_pointer == 83 && y_pointer == 71)
||(x_pointer == 84 && y_pointer == 71)
||(x_pointer == 85 && y_pointer == 71)
||(x_pointer == 86 && y_pointer == 71)
||(x_pointer == 87 && y_pointer == 71)
||(x_pointer == 88 && y_pointer == 71)
||(x_pointer == 89 && y_pointer == 71)
||(x_pointer == 90 && y_pointer == 71)
||(x_pointer == 91 && y_pointer == 71)
||(x_pointer == 92 && y_pointer == 71)
||(x_pointer == 93 && y_pointer == 71)
||(x_pointer == 94 && y_pointer == 71)
||(x_pointer == 95 && y_pointer == 71)
||(x_pointer == 96 && y_pointer == 71)
||(x_pointer == 97 && y_pointer == 71)
||(x_pointer == 98 && y_pointer == 71)
||(x_pointer == 99 && y_pointer == 71)
||(x_pointer == 100 && y_pointer == 71)
||(x_pointer == 101 && y_pointer == 71)
||(x_pointer == 102 && y_pointer == 71)
||(x_pointer == 103 && y_pointer == 71)
||(x_pointer == 104 && y_pointer == 71)
||(x_pointer == 105 && y_pointer == 71)
||(x_pointer == 106 && y_pointer == 71)
||(x_pointer == 107 && y_pointer == 71)
||(x_pointer == 108 && y_pointer == 71)
||(x_pointer == 109 && y_pointer == 71)
||(x_pointer == 110 && y_pointer == 71)
||(x_pointer == 111 && y_pointer == 71)
||(x_pointer == 112 && y_pointer == 71)
||(x_pointer == 113 && y_pointer == 71)
||(x_pointer == 114 && y_pointer == 71)
||(x_pointer == 115 && y_pointer == 71)
||(x_pointer == 50 && y_pointer == 72)
||(x_pointer == 51 && y_pointer == 72)
||(x_pointer == 52 && y_pointer == 72)
||(x_pointer == 53 && y_pointer == 72)
||(x_pointer == 54 && y_pointer == 72)
||(x_pointer == 55 && y_pointer == 72)
||(x_pointer == 56 && y_pointer == 72)
||(x_pointer == 57 && y_pointer == 72)
||(x_pointer == 58 && y_pointer == 72)
||(x_pointer == 59 && y_pointer == 72)
||(x_pointer == 60 && y_pointer == 72)
||(x_pointer == 61 && y_pointer == 72)
||(x_pointer == 62 && y_pointer == 72)
||(x_pointer == 63 && y_pointer == 72)
||(x_pointer == 64 && y_pointer == 72)
||(x_pointer == 65 && y_pointer == 72)
||(x_pointer == 66 && y_pointer == 72)
||(x_pointer == 67 && y_pointer == 72)
||(x_pointer == 68 && y_pointer == 72)
||(x_pointer == 69 && y_pointer == 72)
||(x_pointer == 70 && y_pointer == 72)
||(x_pointer == 71 && y_pointer == 72)
||(x_pointer == 72 && y_pointer == 72)
||(x_pointer == 73 && y_pointer == 72)
||(x_pointer == 74 && y_pointer == 72)
||(x_pointer == 75 && y_pointer == 72)
||(x_pointer == 76 && y_pointer == 72)
||(x_pointer == 77 && y_pointer == 72)
||(x_pointer == 78 && y_pointer == 72)
||(x_pointer == 79 && y_pointer == 72)
||(x_pointer == 80 && y_pointer == 72)
||(x_pointer == 81 && y_pointer == 72)
||(x_pointer == 82 && y_pointer == 72)
||(x_pointer == 83 && y_pointer == 72)
||(x_pointer == 84 && y_pointer == 72)
||(x_pointer == 85 && y_pointer == 72)
||(x_pointer == 86 && y_pointer == 72)
||(x_pointer == 87 && y_pointer == 72)
||(x_pointer == 88 && y_pointer == 72)
||(x_pointer == 89 && y_pointer == 72)
||(x_pointer == 90 && y_pointer == 72)
||(x_pointer == 91 && y_pointer == 72)
||(x_pointer == 92 && y_pointer == 72)
||(x_pointer == 93 && y_pointer == 72)
||(x_pointer == 94 && y_pointer == 72)
||(x_pointer == 95 && y_pointer == 72)
||(x_pointer == 96 && y_pointer == 72)
||(x_pointer == 97 && y_pointer == 72)
||(x_pointer == 98 && y_pointer == 72)
||(x_pointer == 99 && y_pointer == 72)
||(x_pointer == 100 && y_pointer == 72)
||(x_pointer == 101 && y_pointer == 72)
||(x_pointer == 102 && y_pointer == 72)
||(x_pointer == 103 && y_pointer == 72)
||(x_pointer == 104 && y_pointer == 72)
||(x_pointer == 105 && y_pointer == 72)
||(x_pointer == 106 && y_pointer == 72)
||(x_pointer == 107 && y_pointer == 72)
||(x_pointer == 108 && y_pointer == 72)
||(x_pointer == 109 && y_pointer == 72)
||(x_pointer == 110 && y_pointer == 72)
||(x_pointer == 111 && y_pointer == 72)
||(x_pointer == 112 && y_pointer == 72)
||(x_pointer == 113 && y_pointer == 72)
||(x_pointer == 114 && y_pointer == 72)
||(x_pointer == 115 && y_pointer == 72)
||(x_pointer == 50 && y_pointer == 73)
||(x_pointer == 51 && y_pointer == 73)
||(x_pointer == 52 && y_pointer == 73)
||(x_pointer == 53 && y_pointer == 73)
||(x_pointer == 54 && y_pointer == 73)
||(x_pointer == 55 && y_pointer == 73)
||(x_pointer == 56 && y_pointer == 73)
||(x_pointer == 57 && y_pointer == 73)
||(x_pointer == 58 && y_pointer == 73)
||(x_pointer == 59 && y_pointer == 73)
||(x_pointer == 60 && y_pointer == 73)
||(x_pointer == 61 && y_pointer == 73)
||(x_pointer == 62 && y_pointer == 73)
||(x_pointer == 63 && y_pointer == 73)
||(x_pointer == 64 && y_pointer == 73)
||(x_pointer == 65 && y_pointer == 73)
||(x_pointer == 66 && y_pointer == 73)
||(x_pointer == 67 && y_pointer == 73)
||(x_pointer == 68 && y_pointer == 73)
||(x_pointer == 69 && y_pointer == 73)
||(x_pointer == 70 && y_pointer == 73)
||(x_pointer == 71 && y_pointer == 73)
||(x_pointer == 72 && y_pointer == 73)
||(x_pointer == 73 && y_pointer == 73)
||(x_pointer == 74 && y_pointer == 73)
||(x_pointer == 75 && y_pointer == 73)
||(x_pointer == 76 && y_pointer == 73)
||(x_pointer == 77 && y_pointer == 73)
||(x_pointer == 78 && y_pointer == 73)
||(x_pointer == 79 && y_pointer == 73)
||(x_pointer == 80 && y_pointer == 73)
||(x_pointer == 81 && y_pointer == 73)
||(x_pointer == 82 && y_pointer == 73)
||(x_pointer == 83 && y_pointer == 73)
||(x_pointer == 84 && y_pointer == 73)
||(x_pointer == 85 && y_pointer == 73)
||(x_pointer == 86 && y_pointer == 73)
||(x_pointer == 87 && y_pointer == 73)
||(x_pointer == 88 && y_pointer == 73)
||(x_pointer == 89 && y_pointer == 73)
||(x_pointer == 90 && y_pointer == 73)
||(x_pointer == 91 && y_pointer == 73)
||(x_pointer == 92 && y_pointer == 73)
||(x_pointer == 93 && y_pointer == 73)
||(x_pointer == 94 && y_pointer == 73)
||(x_pointer == 95 && y_pointer == 73)
||(x_pointer == 96 && y_pointer == 73)
||(x_pointer == 97 && y_pointer == 73)
||(x_pointer == 98 && y_pointer == 73)
||(x_pointer == 99 && y_pointer == 73)
||(x_pointer == 100 && y_pointer == 73)
||(x_pointer == 101 && y_pointer == 73)
||(x_pointer == 102 && y_pointer == 73)
||(x_pointer == 103 && y_pointer == 73)
||(x_pointer == 104 && y_pointer == 73)
||(x_pointer == 105 && y_pointer == 73)
||(x_pointer == 106 && y_pointer == 73)
||(x_pointer == 107 && y_pointer == 73)
||(x_pointer == 108 && y_pointer == 73)
||(x_pointer == 109 && y_pointer == 73)
||(x_pointer == 110 && y_pointer == 73)
||(x_pointer == 111 && y_pointer == 73)
||(x_pointer == 112 && y_pointer == 73)
||(x_pointer == 113 && y_pointer == 73)
||(x_pointer == 114 && y_pointer == 73)
||(x_pointer == 115 && y_pointer == 73)
||(x_pointer == 50 && y_pointer == 74)
||(x_pointer == 51 && y_pointer == 74)
||(x_pointer == 52 && y_pointer == 74)
||(x_pointer == 53 && y_pointer == 74)
||(x_pointer == 54 && y_pointer == 74)
||(x_pointer == 55 && y_pointer == 74)
||(x_pointer == 56 && y_pointer == 74)
||(x_pointer == 57 && y_pointer == 74)
||(x_pointer == 58 && y_pointer == 74)
||(x_pointer == 59 && y_pointer == 74)
||(x_pointer == 60 && y_pointer == 74)
||(x_pointer == 61 && y_pointer == 74)
||(x_pointer == 62 && y_pointer == 74)
||(x_pointer == 63 && y_pointer == 74)
||(x_pointer == 64 && y_pointer == 74)
||(x_pointer == 65 && y_pointer == 74)
||(x_pointer == 66 && y_pointer == 74)
||(x_pointer == 67 && y_pointer == 74)
||(x_pointer == 68 && y_pointer == 74)
||(x_pointer == 69 && y_pointer == 74)
||(x_pointer == 70 && y_pointer == 74)
||(x_pointer == 71 && y_pointer == 74)
||(x_pointer == 72 && y_pointer == 74)
||(x_pointer == 73 && y_pointer == 74)
||(x_pointer == 74 && y_pointer == 74)
||(x_pointer == 75 && y_pointer == 74)
||(x_pointer == 76 && y_pointer == 74)
||(x_pointer == 77 && y_pointer == 74)
||(x_pointer == 78 && y_pointer == 74)
||(x_pointer == 79 && y_pointer == 74)
||(x_pointer == 80 && y_pointer == 74)
||(x_pointer == 81 && y_pointer == 74)
||(x_pointer == 82 && y_pointer == 74)
||(x_pointer == 83 && y_pointer == 74)
||(x_pointer == 84 && y_pointer == 74)
||(x_pointer == 85 && y_pointer == 74)
||(x_pointer == 86 && y_pointer == 74)
||(x_pointer == 87 && y_pointer == 74)
||(x_pointer == 88 && y_pointer == 74)
||(x_pointer == 89 && y_pointer == 74)
||(x_pointer == 90 && y_pointer == 74)
||(x_pointer == 91 && y_pointer == 74)
||(x_pointer == 92 && y_pointer == 74)
||(x_pointer == 93 && y_pointer == 74)
||(x_pointer == 94 && y_pointer == 74)
||(x_pointer == 95 && y_pointer == 74)
||(x_pointer == 96 && y_pointer == 74)
||(x_pointer == 97 && y_pointer == 74)
||(x_pointer == 98 && y_pointer == 74)
||(x_pointer == 99 && y_pointer == 74)
||(x_pointer == 100 && y_pointer == 74)
||(x_pointer == 101 && y_pointer == 74)
||(x_pointer == 102 && y_pointer == 74)
||(x_pointer == 103 && y_pointer == 74)
||(x_pointer == 104 && y_pointer == 74)
||(x_pointer == 105 && y_pointer == 74)
||(x_pointer == 106 && y_pointer == 74)
||(x_pointer == 107 && y_pointer == 74)
||(x_pointer == 108 && y_pointer == 74)
||(x_pointer == 109 && y_pointer == 74)
||(x_pointer == 110 && y_pointer == 74)
||(x_pointer == 111 && y_pointer == 74)
||(x_pointer == 112 && y_pointer == 74)
||(x_pointer == 113 && y_pointer == 74)
||(x_pointer == 114 && y_pointer == 74)
||(x_pointer == 115 && y_pointer == 74)
||(x_pointer == 50 && y_pointer == 75)
||(x_pointer == 51 && y_pointer == 75)
||(x_pointer == 52 && y_pointer == 75)
||(x_pointer == 53 && y_pointer == 75)
||(x_pointer == 54 && y_pointer == 75)
||(x_pointer == 55 && y_pointer == 75)
||(x_pointer == 56 && y_pointer == 75)
||(x_pointer == 57 && y_pointer == 75)
||(x_pointer == 58 && y_pointer == 75)
||(x_pointer == 59 && y_pointer == 75)
||(x_pointer == 60 && y_pointer == 75)
||(x_pointer == 61 && y_pointer == 75)
||(x_pointer == 62 && y_pointer == 75)
||(x_pointer == 63 && y_pointer == 75)
||(x_pointer == 64 && y_pointer == 75)
||(x_pointer == 65 && y_pointer == 75)
||(x_pointer == 66 && y_pointer == 75)
||(x_pointer == 67 && y_pointer == 75)
||(x_pointer == 68 && y_pointer == 75)
||(x_pointer == 69 && y_pointer == 75)
||(x_pointer == 70 && y_pointer == 75)
||(x_pointer == 71 && y_pointer == 75)
||(x_pointer == 72 && y_pointer == 75)
||(x_pointer == 73 && y_pointer == 75)
||(x_pointer == 74 && y_pointer == 75)
||(x_pointer == 75 && y_pointer == 75)
||(x_pointer == 76 && y_pointer == 75)
||(x_pointer == 77 && y_pointer == 75)
||(x_pointer == 78 && y_pointer == 75)
||(x_pointer == 79 && y_pointer == 75)
||(x_pointer == 80 && y_pointer == 75)
||(x_pointer == 81 && y_pointer == 75)
||(x_pointer == 82 && y_pointer == 75)
||(x_pointer == 83 && y_pointer == 75)
||(x_pointer == 84 && y_pointer == 75)
||(x_pointer == 85 && y_pointer == 75)
||(x_pointer == 86 && y_pointer == 75)
||(x_pointer == 87 && y_pointer == 75)
||(x_pointer == 88 && y_pointer == 75)
||(x_pointer == 89 && y_pointer == 75)
||(x_pointer == 90 && y_pointer == 75)
||(x_pointer == 91 && y_pointer == 75)
||(x_pointer == 92 && y_pointer == 75)
||(x_pointer == 93 && y_pointer == 75)
||(x_pointer == 94 && y_pointer == 75)
||(x_pointer == 95 && y_pointer == 75)
||(x_pointer == 96 && y_pointer == 75)
||(x_pointer == 97 && y_pointer == 75)
||(x_pointer == 98 && y_pointer == 75)
||(x_pointer == 99 && y_pointer == 75)
||(x_pointer == 100 && y_pointer == 75)
||(x_pointer == 101 && y_pointer == 75)
||(x_pointer == 102 && y_pointer == 75)
||(x_pointer == 103 && y_pointer == 75)
||(x_pointer == 104 && y_pointer == 75)
||(x_pointer == 105 && y_pointer == 75)
||(x_pointer == 106 && y_pointer == 75)
||(x_pointer == 107 && y_pointer == 75)
||(x_pointer == 108 && y_pointer == 75)
||(x_pointer == 109 && y_pointer == 75)
||(x_pointer == 110 && y_pointer == 75)
||(x_pointer == 111 && y_pointer == 75)
||(x_pointer == 112 && y_pointer == 75)
||(x_pointer == 113 && y_pointer == 75)
||(x_pointer == 114 && y_pointer == 75)
||(x_pointer == 115 && y_pointer == 75)
||(x_pointer == 50 && y_pointer == 76)
||(x_pointer == 51 && y_pointer == 76)
||(x_pointer == 52 && y_pointer == 76)
||(x_pointer == 53 && y_pointer == 76)
||(x_pointer == 54 && y_pointer == 76)
||(x_pointer == 55 && y_pointer == 76)
||(x_pointer == 56 && y_pointer == 76)
||(x_pointer == 57 && y_pointer == 76)
||(x_pointer == 58 && y_pointer == 76)
||(x_pointer == 59 && y_pointer == 76)
||(x_pointer == 60 && y_pointer == 76)
||(x_pointer == 61 && y_pointer == 76)
||(x_pointer == 62 && y_pointer == 76)
||(x_pointer == 63 && y_pointer == 76)
||(x_pointer == 64 && y_pointer == 76)
||(x_pointer == 65 && y_pointer == 76)
||(x_pointer == 66 && y_pointer == 76)
||(x_pointer == 67 && y_pointer == 76)
||(x_pointer == 68 && y_pointer == 76)
||(x_pointer == 69 && y_pointer == 76)
||(x_pointer == 70 && y_pointer == 76)
||(x_pointer == 71 && y_pointer == 76)
||(x_pointer == 72 && y_pointer == 76)
||(x_pointer == 73 && y_pointer == 76)
||(x_pointer == 74 && y_pointer == 76)
||(x_pointer == 75 && y_pointer == 76)
||(x_pointer == 76 && y_pointer == 76)
||(x_pointer == 77 && y_pointer == 76)
||(x_pointer == 78 && y_pointer == 76)
||(x_pointer == 79 && y_pointer == 76)
||(x_pointer == 80 && y_pointer == 76)
||(x_pointer == 81 && y_pointer == 76)
||(x_pointer == 82 && y_pointer == 76)
||(x_pointer == 83 && y_pointer == 76)
||(x_pointer == 84 && y_pointer == 76)
||(x_pointer == 85 && y_pointer == 76)
||(x_pointer == 86 && y_pointer == 76)
||(x_pointer == 87 && y_pointer == 76)
||(x_pointer == 88 && y_pointer == 76)
||(x_pointer == 89 && y_pointer == 76)
||(x_pointer == 90 && y_pointer == 76)
||(x_pointer == 91 && y_pointer == 76)
||(x_pointer == 92 && y_pointer == 76)
||(x_pointer == 93 && y_pointer == 76)
||(x_pointer == 94 && y_pointer == 76)
||(x_pointer == 95 && y_pointer == 76)
||(x_pointer == 96 && y_pointer == 76)
||(x_pointer == 97 && y_pointer == 76)
||(x_pointer == 98 && y_pointer == 76)
||(x_pointer == 99 && y_pointer == 76)
||(x_pointer == 100 && y_pointer == 76)
||(x_pointer == 101 && y_pointer == 76)
||(x_pointer == 102 && y_pointer == 76)
||(x_pointer == 103 && y_pointer == 76)
||(x_pointer == 104 && y_pointer == 76)
||(x_pointer == 105 && y_pointer == 76)
||(x_pointer == 106 && y_pointer == 76)
||(x_pointer == 107 && y_pointer == 76)
||(x_pointer == 108 && y_pointer == 76)
||(x_pointer == 109 && y_pointer == 76)
||(x_pointer == 110 && y_pointer == 76)
||(x_pointer == 111 && y_pointer == 76)
||(x_pointer == 112 && y_pointer == 76)
||(x_pointer == 113 && y_pointer == 76)
||(x_pointer == 114 && y_pointer == 76)
||(x_pointer == 115 && y_pointer == 76)
||(x_pointer == 23 && y_pointer == 79)
||(x_pointer == 24 && y_pointer == 79)
||(x_pointer == 25 && y_pointer == 79)
||(x_pointer == 26 && y_pointer == 79)
||(x_pointer == 27 && y_pointer == 79)
||(x_pointer == 28 && y_pointer == 79)
||(x_pointer == 29 && y_pointer == 79)
||(x_pointer == 30 && y_pointer == 79)
||(x_pointer == 31 && y_pointer == 79)
||(x_pointer == 23 && y_pointer == 80)
||(x_pointer == 24 && y_pointer == 80)
||(x_pointer == 25 && y_pointer == 80)
||(x_pointer == 26 && y_pointer == 80)
||(x_pointer == 27 && y_pointer == 80)
||(x_pointer == 28 && y_pointer == 80)
||(x_pointer == 29 && y_pointer == 80)
||(x_pointer == 30 && y_pointer == 80)
||(x_pointer == 31 && y_pointer == 80)
||(x_pointer == 134 && y_pointer == 80)
||(x_pointer == 135 && y_pointer == 80)
||(x_pointer == 136 && y_pointer == 80)
||(x_pointer == 137 && y_pointer == 80)
||(x_pointer == 138 && y_pointer == 80)
||(x_pointer == 139 && y_pointer == 80)
||(x_pointer == 140 && y_pointer == 80)
||(x_pointer == 141 && y_pointer == 80)
||(x_pointer == 142 && y_pointer == 80)
||(x_pointer == 23 && y_pointer == 81)
||(x_pointer == 24 && y_pointer == 81)
||(x_pointer == 25 && y_pointer == 81)
||(x_pointer == 26 && y_pointer == 81)
||(x_pointer == 27 && y_pointer == 81)
||(x_pointer == 28 && y_pointer == 81)
||(x_pointer == 29 && y_pointer == 81)
||(x_pointer == 30 && y_pointer == 81)
||(x_pointer == 31 && y_pointer == 81)
||(x_pointer == 134 && y_pointer == 81)
||(x_pointer == 135 && y_pointer == 81)
||(x_pointer == 136 && y_pointer == 81)
||(x_pointer == 137 && y_pointer == 81)
||(x_pointer == 138 && y_pointer == 81)
||(x_pointer == 139 && y_pointer == 81)
||(x_pointer == 140 && y_pointer == 81)
||(x_pointer == 141 && y_pointer == 81)
||(x_pointer == 142 && y_pointer == 81)
||(x_pointer == 23 && y_pointer == 82)
||(x_pointer == 24 && y_pointer == 82)
||(x_pointer == 25 && y_pointer == 82)
||(x_pointer == 26 && y_pointer == 82)
||(x_pointer == 27 && y_pointer == 82)
||(x_pointer == 28 && y_pointer == 82)
||(x_pointer == 29 && y_pointer == 82)
||(x_pointer == 30 && y_pointer == 82)
||(x_pointer == 31 && y_pointer == 82)
||(x_pointer == 134 && y_pointer == 82)
||(x_pointer == 135 && y_pointer == 82)
||(x_pointer == 136 && y_pointer == 82)
||(x_pointer == 137 && y_pointer == 82)
||(x_pointer == 138 && y_pointer == 82)
||(x_pointer == 139 && y_pointer == 82)
||(x_pointer == 140 && y_pointer == 82)
||(x_pointer == 141 && y_pointer == 82)
||(x_pointer == 142 && y_pointer == 82)
||(x_pointer == 23 && y_pointer == 83)
||(x_pointer == 24 && y_pointer == 83)
||(x_pointer == 25 && y_pointer == 83)
||(x_pointer == 26 && y_pointer == 83)
||(x_pointer == 27 && y_pointer == 83)
||(x_pointer == 28 && y_pointer == 83)
||(x_pointer == 29 && y_pointer == 83)
||(x_pointer == 30 && y_pointer == 83)
||(x_pointer == 31 && y_pointer == 83)
||(x_pointer == 134 && y_pointer == 83)
||(x_pointer == 135 && y_pointer == 83)
||(x_pointer == 136 && y_pointer == 83)
||(x_pointer == 137 && y_pointer == 83)
||(x_pointer == 138 && y_pointer == 83)
||(x_pointer == 139 && y_pointer == 83)
||(x_pointer == 140 && y_pointer == 83)
||(x_pointer == 141 && y_pointer == 83)
||(x_pointer == 142 && y_pointer == 83)
||(x_pointer == 23 && y_pointer == 84)
||(x_pointer == 24 && y_pointer == 84)
||(x_pointer == 25 && y_pointer == 84)
||(x_pointer == 26 && y_pointer == 84)
||(x_pointer == 27 && y_pointer == 84)
||(x_pointer == 28 && y_pointer == 84)
||(x_pointer == 29 && y_pointer == 84)
||(x_pointer == 30 && y_pointer == 84)
||(x_pointer == 31 && y_pointer == 84)
||(x_pointer == 134 && y_pointer == 84)
||(x_pointer == 135 && y_pointer == 84)
||(x_pointer == 136 && y_pointer == 84)
||(x_pointer == 137 && y_pointer == 84)
||(x_pointer == 138 && y_pointer == 84)
||(x_pointer == 139 && y_pointer == 84)
||(x_pointer == 140 && y_pointer == 84)
||(x_pointer == 141 && y_pointer == 84)
||(x_pointer == 142 && y_pointer == 84)
||(x_pointer == 23 && y_pointer == 85)
||(x_pointer == 24 && y_pointer == 85)
||(x_pointer == 25 && y_pointer == 85)
||(x_pointer == 26 && y_pointer == 85)
||(x_pointer == 27 && y_pointer == 85)
||(x_pointer == 28 && y_pointer == 85)
||(x_pointer == 29 && y_pointer == 85)
||(x_pointer == 30 && y_pointer == 85)
||(x_pointer == 31 && y_pointer == 85)
||(x_pointer == 134 && y_pointer == 85)
||(x_pointer == 135 && y_pointer == 85)
||(x_pointer == 136 && y_pointer == 85)
||(x_pointer == 137 && y_pointer == 85)
||(x_pointer == 138 && y_pointer == 85)
||(x_pointer == 139 && y_pointer == 85)
||(x_pointer == 140 && y_pointer == 85)
||(x_pointer == 141 && y_pointer == 85)
||(x_pointer == 142 && y_pointer == 85)
||(x_pointer == 23 && y_pointer == 86)
||(x_pointer == 24 && y_pointer == 86)
||(x_pointer == 25 && y_pointer == 86)
||(x_pointer == 26 && y_pointer == 86)
||(x_pointer == 27 && y_pointer == 86)
||(x_pointer == 28 && y_pointer == 86)
||(x_pointer == 29 && y_pointer == 86)
||(x_pointer == 30 && y_pointer == 86)
||(x_pointer == 31 && y_pointer == 86)
||(x_pointer == 134 && y_pointer == 86)
||(x_pointer == 135 && y_pointer == 86)
||(x_pointer == 136 && y_pointer == 86)
||(x_pointer == 137 && y_pointer == 86)
||(x_pointer == 138 && y_pointer == 86)
||(x_pointer == 139 && y_pointer == 86)
||(x_pointer == 140 && y_pointer == 86)
||(x_pointer == 141 && y_pointer == 86)
||(x_pointer == 142 && y_pointer == 86)
||(x_pointer == 23 && y_pointer == 87)
||(x_pointer == 24 && y_pointer == 87)
||(x_pointer == 25 && y_pointer == 87)
||(x_pointer == 26 && y_pointer == 87)
||(x_pointer == 27 && y_pointer == 87)
||(x_pointer == 28 && y_pointer == 87)
||(x_pointer == 29 && y_pointer == 87)
||(x_pointer == 30 && y_pointer == 87)
||(x_pointer == 31 && y_pointer == 87)
||(x_pointer == 134 && y_pointer == 87)
||(x_pointer == 135 && y_pointer == 87)
||(x_pointer == 136 && y_pointer == 87)
||(x_pointer == 137 && y_pointer == 87)
||(x_pointer == 138 && y_pointer == 87)
||(x_pointer == 139 && y_pointer == 87)
||(x_pointer == 140 && y_pointer == 87)
||(x_pointer == 141 && y_pointer == 87)
||(x_pointer == 142 && y_pointer == 87)
||(x_pointer == 23 && y_pointer == 88)
||(x_pointer == 24 && y_pointer == 88)
||(x_pointer == 25 && y_pointer == 88)
||(x_pointer == 26 && y_pointer == 88)
||(x_pointer == 27 && y_pointer == 88)
||(x_pointer == 28 && y_pointer == 88)
||(x_pointer == 29 && y_pointer == 88)
||(x_pointer == 30 && y_pointer == 88)
||(x_pointer == 31 && y_pointer == 88)
||(x_pointer == 134 && y_pointer == 88)
||(x_pointer == 135 && y_pointer == 88)
||(x_pointer == 136 && y_pointer == 88)
||(x_pointer == 137 && y_pointer == 88)
||(x_pointer == 138 && y_pointer == 88)
||(x_pointer == 139 && y_pointer == 88)
||(x_pointer == 140 && y_pointer == 88)
||(x_pointer == 141 && y_pointer == 88)
||(x_pointer == 142 && y_pointer == 88)
||(x_pointer == 23 && y_pointer == 89)
||(x_pointer == 24 && y_pointer == 89)
||(x_pointer == 25 && y_pointer == 89)
||(x_pointer == 26 && y_pointer == 89)
||(x_pointer == 27 && y_pointer == 89)
||(x_pointer == 28 && y_pointer == 89)
||(x_pointer == 29 && y_pointer == 89)
||(x_pointer == 30 && y_pointer == 89)
||(x_pointer == 31 && y_pointer == 89)
||(x_pointer == 134 && y_pointer == 89)
||(x_pointer == 135 && y_pointer == 89)
||(x_pointer == 136 && y_pointer == 89)
||(x_pointer == 137 && y_pointer == 89)
||(x_pointer == 138 && y_pointer == 89)
||(x_pointer == 139 && y_pointer == 89)
||(x_pointer == 140 && y_pointer == 89)
||(x_pointer == 141 && y_pointer == 89)
||(x_pointer == 142 && y_pointer == 89)
||(x_pointer == 23 && y_pointer == 90)
||(x_pointer == 24 && y_pointer == 90)
||(x_pointer == 25 && y_pointer == 90)
||(x_pointer == 26 && y_pointer == 90)
||(x_pointer == 27 && y_pointer == 90)
||(x_pointer == 28 && y_pointer == 90)
||(x_pointer == 29 && y_pointer == 90)
||(x_pointer == 30 && y_pointer == 90)
||(x_pointer == 31 && y_pointer == 90)
||(x_pointer == 134 && y_pointer == 90)
||(x_pointer == 135 && y_pointer == 90)
||(x_pointer == 136 && y_pointer == 90)
||(x_pointer == 137 && y_pointer == 90)
||(x_pointer == 138 && y_pointer == 90)
||(x_pointer == 139 && y_pointer == 90)
||(x_pointer == 140 && y_pointer == 90)
||(x_pointer == 141 && y_pointer == 90)
||(x_pointer == 142 && y_pointer == 90)
||(x_pointer == 23 && y_pointer == 91)
||(x_pointer == 24 && y_pointer == 91)
||(x_pointer == 25 && y_pointer == 91)
||(x_pointer == 26 && y_pointer == 91)
||(x_pointer == 27 && y_pointer == 91)
||(x_pointer == 28 && y_pointer == 91)
||(x_pointer == 29 && y_pointer == 91)
||(x_pointer == 30 && y_pointer == 91)
||(x_pointer == 31 && y_pointer == 91)
||(x_pointer == 134 && y_pointer == 91)
||(x_pointer == 135 && y_pointer == 91)
||(x_pointer == 136 && y_pointer == 91)
||(x_pointer == 137 && y_pointer == 91)
||(x_pointer == 138 && y_pointer == 91)
||(x_pointer == 139 && y_pointer == 91)
||(x_pointer == 140 && y_pointer == 91)
||(x_pointer == 141 && y_pointer == 91)
||(x_pointer == 142 && y_pointer == 91)
||(x_pointer == 23 && y_pointer == 92)
||(x_pointer == 24 && y_pointer == 92)
||(x_pointer == 25 && y_pointer == 92)
||(x_pointer == 26 && y_pointer == 92)
||(x_pointer == 27 && y_pointer == 92)
||(x_pointer == 28 && y_pointer == 92)
||(x_pointer == 29 && y_pointer == 92)
||(x_pointer == 30 && y_pointer == 92)
||(x_pointer == 31 && y_pointer == 92)
||(x_pointer == 122 && y_pointer == 92)
||(x_pointer == 123 && y_pointer == 92)
||(x_pointer == 124 && y_pointer == 92)
||(x_pointer == 125 && y_pointer == 92)
||(x_pointer == 126 && y_pointer == 92)
||(x_pointer == 127 && y_pointer == 92)
||(x_pointer == 128 && y_pointer == 92)
||(x_pointer == 129 && y_pointer == 92)
||(x_pointer == 130 && y_pointer == 92)
||(x_pointer == 131 && y_pointer == 92)
||(x_pointer == 132 && y_pointer == 92)
||(x_pointer == 133 && y_pointer == 92)
||(x_pointer == 134 && y_pointer == 92)
||(x_pointer == 135 && y_pointer == 92)
||(x_pointer == 136 && y_pointer == 92)
||(x_pointer == 137 && y_pointer == 92)
||(x_pointer == 138 && y_pointer == 92)
||(x_pointer == 139 && y_pointer == 92)
||(x_pointer == 140 && y_pointer == 92)
||(x_pointer == 141 && y_pointer == 92)
||(x_pointer == 142 && y_pointer == 92)
||(x_pointer == 23 && y_pointer == 93)
||(x_pointer == 24 && y_pointer == 93)
||(x_pointer == 25 && y_pointer == 93)
||(x_pointer == 26 && y_pointer == 93)
||(x_pointer == 27 && y_pointer == 93)
||(x_pointer == 28 && y_pointer == 93)
||(x_pointer == 29 && y_pointer == 93)
||(x_pointer == 30 && y_pointer == 93)
||(x_pointer == 31 && y_pointer == 93)
||(x_pointer == 32 && y_pointer == 93)
||(x_pointer == 33 && y_pointer == 93)
||(x_pointer == 34 && y_pointer == 93)
||(x_pointer == 35 && y_pointer == 93)
||(x_pointer == 36 && y_pointer == 93)
||(x_pointer == 37 && y_pointer == 93)
||(x_pointer == 38 && y_pointer == 93)
||(x_pointer == 39 && y_pointer == 93)
||(x_pointer == 40 && y_pointer == 93)
||(x_pointer == 41 && y_pointer == 93)
||(x_pointer == 42 && y_pointer == 93)
||(x_pointer == 43 && y_pointer == 93)
||(x_pointer == 122 && y_pointer == 93)
||(x_pointer == 123 && y_pointer == 93)
||(x_pointer == 124 && y_pointer == 93)
||(x_pointer == 125 && y_pointer == 93)
||(x_pointer == 126 && y_pointer == 93)
||(x_pointer == 127 && y_pointer == 93)
||(x_pointer == 128 && y_pointer == 93)
||(x_pointer == 129 && y_pointer == 93)
||(x_pointer == 130 && y_pointer == 93)
||(x_pointer == 131 && y_pointer == 93)
||(x_pointer == 132 && y_pointer == 93)
||(x_pointer == 133 && y_pointer == 93)
||(x_pointer == 134 && y_pointer == 93)
||(x_pointer == 135 && y_pointer == 93)
||(x_pointer == 136 && y_pointer == 93)
||(x_pointer == 137 && y_pointer == 93)
||(x_pointer == 138 && y_pointer == 93)
||(x_pointer == 139 && y_pointer == 93)
||(x_pointer == 140 && y_pointer == 93)
||(x_pointer == 141 && y_pointer == 93)
||(x_pointer == 142 && y_pointer == 93)
||(x_pointer == 23 && y_pointer == 94)
||(x_pointer == 24 && y_pointer == 94)
||(x_pointer == 25 && y_pointer == 94)
||(x_pointer == 26 && y_pointer == 94)
||(x_pointer == 27 && y_pointer == 94)
||(x_pointer == 28 && y_pointer == 94)
||(x_pointer == 29 && y_pointer == 94)
||(x_pointer == 30 && y_pointer == 94)
||(x_pointer == 31 && y_pointer == 94)
||(x_pointer == 32 && y_pointer == 94)
||(x_pointer == 33 && y_pointer == 94)
||(x_pointer == 34 && y_pointer == 94)
||(x_pointer == 35 && y_pointer == 94)
||(x_pointer == 36 && y_pointer == 94)
||(x_pointer == 37 && y_pointer == 94)
||(x_pointer == 38 && y_pointer == 94)
||(x_pointer == 39 && y_pointer == 94)
||(x_pointer == 40 && y_pointer == 94)
||(x_pointer == 41 && y_pointer == 94)
||(x_pointer == 42 && y_pointer == 94)
||(x_pointer == 43 && y_pointer == 94)
||(x_pointer == 122 && y_pointer == 94)
||(x_pointer == 123 && y_pointer == 94)
||(x_pointer == 124 && y_pointer == 94)
||(x_pointer == 125 && y_pointer == 94)
||(x_pointer == 126 && y_pointer == 94)
||(x_pointer == 127 && y_pointer == 94)
||(x_pointer == 128 && y_pointer == 94)
||(x_pointer == 129 && y_pointer == 94)
||(x_pointer == 130 && y_pointer == 94)
||(x_pointer == 131 && y_pointer == 94)
||(x_pointer == 132 && y_pointer == 94)
||(x_pointer == 133 && y_pointer == 94)
||(x_pointer == 134 && y_pointer == 94)
||(x_pointer == 135 && y_pointer == 94)
||(x_pointer == 136 && y_pointer == 94)
||(x_pointer == 137 && y_pointer == 94)
||(x_pointer == 138 && y_pointer == 94)
||(x_pointer == 139 && y_pointer == 94)
||(x_pointer == 140 && y_pointer == 94)
||(x_pointer == 141 && y_pointer == 94)
||(x_pointer == 142 && y_pointer == 94)
||(x_pointer == 23 && y_pointer == 95)
||(x_pointer == 24 && y_pointer == 95)
||(x_pointer == 25 && y_pointer == 95)
||(x_pointer == 26 && y_pointer == 95)
||(x_pointer == 27 && y_pointer == 95)
||(x_pointer == 28 && y_pointer == 95)
||(x_pointer == 29 && y_pointer == 95)
||(x_pointer == 30 && y_pointer == 95)
||(x_pointer == 31 && y_pointer == 95)
||(x_pointer == 32 && y_pointer == 95)
||(x_pointer == 33 && y_pointer == 95)
||(x_pointer == 34 && y_pointer == 95)
||(x_pointer == 35 && y_pointer == 95)
||(x_pointer == 36 && y_pointer == 95)
||(x_pointer == 37 && y_pointer == 95)
||(x_pointer == 38 && y_pointer == 95)
||(x_pointer == 39 && y_pointer == 95)
||(x_pointer == 40 && y_pointer == 95)
||(x_pointer == 41 && y_pointer == 95)
||(x_pointer == 42 && y_pointer == 95)
||(x_pointer == 43 && y_pointer == 95)
||(x_pointer == 122 && y_pointer == 95)
||(x_pointer == 123 && y_pointer == 95)
||(x_pointer == 124 && y_pointer == 95)
||(x_pointer == 125 && y_pointer == 95)
||(x_pointer == 126 && y_pointer == 95)
||(x_pointer == 127 && y_pointer == 95)
||(x_pointer == 128 && y_pointer == 95)
||(x_pointer == 129 && y_pointer == 95)
||(x_pointer == 130 && y_pointer == 95)
||(x_pointer == 131 && y_pointer == 95)
||(x_pointer == 132 && y_pointer == 95)
||(x_pointer == 133 && y_pointer == 95)
||(x_pointer == 134 && y_pointer == 95)
||(x_pointer == 135 && y_pointer == 95)
||(x_pointer == 136 && y_pointer == 95)
||(x_pointer == 137 && y_pointer == 95)
||(x_pointer == 138 && y_pointer == 95)
||(x_pointer == 139 && y_pointer == 95)
||(x_pointer == 140 && y_pointer == 95)
||(x_pointer == 141 && y_pointer == 95)
||(x_pointer == 142 && y_pointer == 95)
||(x_pointer == 23 && y_pointer == 96)
||(x_pointer == 24 && y_pointer == 96)
||(x_pointer == 25 && y_pointer == 96)
||(x_pointer == 26 && y_pointer == 96)
||(x_pointer == 27 && y_pointer == 96)
||(x_pointer == 28 && y_pointer == 96)
||(x_pointer == 29 && y_pointer == 96)
||(x_pointer == 30 && y_pointer == 96)
||(x_pointer == 31 && y_pointer == 96)
||(x_pointer == 32 && y_pointer == 96)
||(x_pointer == 33 && y_pointer == 96)
||(x_pointer == 34 && y_pointer == 96)
||(x_pointer == 35 && y_pointer == 96)
||(x_pointer == 36 && y_pointer == 96)
||(x_pointer == 37 && y_pointer == 96)
||(x_pointer == 38 && y_pointer == 96)
||(x_pointer == 39 && y_pointer == 96)
||(x_pointer == 40 && y_pointer == 96)
||(x_pointer == 41 && y_pointer == 96)
||(x_pointer == 42 && y_pointer == 96)
||(x_pointer == 43 && y_pointer == 96)
||(x_pointer == 122 && y_pointer == 96)
||(x_pointer == 123 && y_pointer == 96)
||(x_pointer == 124 && y_pointer == 96)
||(x_pointer == 125 && y_pointer == 96)
||(x_pointer == 126 && y_pointer == 96)
||(x_pointer == 127 && y_pointer == 96)
||(x_pointer == 128 && y_pointer == 96)
||(x_pointer == 129 && y_pointer == 96)
||(x_pointer == 130 && y_pointer == 96)
||(x_pointer == 131 && y_pointer == 96)
||(x_pointer == 132 && y_pointer == 96)
||(x_pointer == 133 && y_pointer == 96)
||(x_pointer == 134 && y_pointer == 96)
||(x_pointer == 135 && y_pointer == 96)
||(x_pointer == 136 && y_pointer == 96)
||(x_pointer == 137 && y_pointer == 96)
||(x_pointer == 138 && y_pointer == 96)
||(x_pointer == 139 && y_pointer == 96)
||(x_pointer == 140 && y_pointer == 96)
||(x_pointer == 141 && y_pointer == 96)
||(x_pointer == 142 && y_pointer == 96)
||(x_pointer == 23 && y_pointer == 97)
||(x_pointer == 24 && y_pointer == 97)
||(x_pointer == 25 && y_pointer == 97)
||(x_pointer == 26 && y_pointer == 97)
||(x_pointer == 27 && y_pointer == 97)
||(x_pointer == 28 && y_pointer == 97)
||(x_pointer == 29 && y_pointer == 97)
||(x_pointer == 30 && y_pointer == 97)
||(x_pointer == 31 && y_pointer == 97)
||(x_pointer == 32 && y_pointer == 97)
||(x_pointer == 33 && y_pointer == 97)
||(x_pointer == 34 && y_pointer == 97)
||(x_pointer == 35 && y_pointer == 97)
||(x_pointer == 36 && y_pointer == 97)
||(x_pointer == 37 && y_pointer == 97)
||(x_pointer == 38 && y_pointer == 97)
||(x_pointer == 39 && y_pointer == 97)
||(x_pointer == 40 && y_pointer == 97)
||(x_pointer == 41 && y_pointer == 97)
||(x_pointer == 42 && y_pointer == 97)
||(x_pointer == 43 && y_pointer == 97)
||(x_pointer == 122 && y_pointer == 97)
||(x_pointer == 123 && y_pointer == 97)
||(x_pointer == 124 && y_pointer == 97)
||(x_pointer == 125 && y_pointer == 97)
||(x_pointer == 126 && y_pointer == 97)
||(x_pointer == 127 && y_pointer == 97)
||(x_pointer == 128 && y_pointer == 97)
||(x_pointer == 129 && y_pointer == 97)
||(x_pointer == 130 && y_pointer == 97)
||(x_pointer == 131 && y_pointer == 97)
||(x_pointer == 132 && y_pointer == 97)
||(x_pointer == 133 && y_pointer == 97)
||(x_pointer == 134 && y_pointer == 97)
||(x_pointer == 135 && y_pointer == 97)
||(x_pointer == 136 && y_pointer == 97)
||(x_pointer == 137 && y_pointer == 97)
||(x_pointer == 138 && y_pointer == 97)
||(x_pointer == 139 && y_pointer == 97)
||(x_pointer == 140 && y_pointer == 97)
||(x_pointer == 141 && y_pointer == 97)
||(x_pointer == 142 && y_pointer == 97)
||(x_pointer == 23 && y_pointer == 98)
||(x_pointer == 24 && y_pointer == 98)
||(x_pointer == 25 && y_pointer == 98)
||(x_pointer == 26 && y_pointer == 98)
||(x_pointer == 27 && y_pointer == 98)
||(x_pointer == 28 && y_pointer == 98)
||(x_pointer == 29 && y_pointer == 98)
||(x_pointer == 30 && y_pointer == 98)
||(x_pointer == 31 && y_pointer == 98)
||(x_pointer == 32 && y_pointer == 98)
||(x_pointer == 33 && y_pointer == 98)
||(x_pointer == 34 && y_pointer == 98)
||(x_pointer == 35 && y_pointer == 98)
||(x_pointer == 36 && y_pointer == 98)
||(x_pointer == 37 && y_pointer == 98)
||(x_pointer == 38 && y_pointer == 98)
||(x_pointer == 39 && y_pointer == 98)
||(x_pointer == 40 && y_pointer == 98)
||(x_pointer == 41 && y_pointer == 98)
||(x_pointer == 42 && y_pointer == 98)
||(x_pointer == 43 && y_pointer == 98)
||(x_pointer == 122 && y_pointer == 98)
||(x_pointer == 123 && y_pointer == 98)
||(x_pointer == 124 && y_pointer == 98)
||(x_pointer == 125 && y_pointer == 98)
||(x_pointer == 126 && y_pointer == 98)
||(x_pointer == 127 && y_pointer == 98)
||(x_pointer == 128 && y_pointer == 98)
||(x_pointer == 129 && y_pointer == 98)
||(x_pointer == 130 && y_pointer == 98)
||(x_pointer == 131 && y_pointer == 98)
||(x_pointer == 132 && y_pointer == 98)
||(x_pointer == 133 && y_pointer == 98)
||(x_pointer == 134 && y_pointer == 98)
||(x_pointer == 135 && y_pointer == 98)
||(x_pointer == 136 && y_pointer == 98)
||(x_pointer == 137 && y_pointer == 98)
||(x_pointer == 138 && y_pointer == 98)
||(x_pointer == 139 && y_pointer == 98)
||(x_pointer == 140 && y_pointer == 98)
||(x_pointer == 141 && y_pointer == 98)
||(x_pointer == 142 && y_pointer == 98)
||(x_pointer == 23 && y_pointer == 99)
||(x_pointer == 24 && y_pointer == 99)
||(x_pointer == 25 && y_pointer == 99)
||(x_pointer == 26 && y_pointer == 99)
||(x_pointer == 27 && y_pointer == 99)
||(x_pointer == 28 && y_pointer == 99)
||(x_pointer == 29 && y_pointer == 99)
||(x_pointer == 30 && y_pointer == 99)
||(x_pointer == 31 && y_pointer == 99)
||(x_pointer == 32 && y_pointer == 99)
||(x_pointer == 33 && y_pointer == 99)
||(x_pointer == 34 && y_pointer == 99)
||(x_pointer == 35 && y_pointer == 99)
||(x_pointer == 36 && y_pointer == 99)
||(x_pointer == 37 && y_pointer == 99)
||(x_pointer == 38 && y_pointer == 99)
||(x_pointer == 39 && y_pointer == 99)
||(x_pointer == 40 && y_pointer == 99)
||(x_pointer == 41 && y_pointer == 99)
||(x_pointer == 42 && y_pointer == 99)
||(x_pointer == 43 && y_pointer == 99)
||(x_pointer == 122 && y_pointer == 99)
||(x_pointer == 123 && y_pointer == 99)
||(x_pointer == 124 && y_pointer == 99)
||(x_pointer == 125 && y_pointer == 99)
||(x_pointer == 126 && y_pointer == 99)
||(x_pointer == 127 && y_pointer == 99)
||(x_pointer == 128 && y_pointer == 99)
||(x_pointer == 129 && y_pointer == 99)
||(x_pointer == 130 && y_pointer == 99)
||(x_pointer == 131 && y_pointer == 99)
||(x_pointer == 132 && y_pointer == 99)
||(x_pointer == 133 && y_pointer == 99)
||(x_pointer == 134 && y_pointer == 99)
||(x_pointer == 135 && y_pointer == 99)
||(x_pointer == 136 && y_pointer == 99)
||(x_pointer == 137 && y_pointer == 99)
||(x_pointer == 138 && y_pointer == 99)
||(x_pointer == 139 && y_pointer == 99)
||(x_pointer == 140 && y_pointer == 99)
||(x_pointer == 141 && y_pointer == 99)
||(x_pointer == 142 && y_pointer == 99)
||(x_pointer == 23 && y_pointer == 100)
||(x_pointer == 24 && y_pointer == 100)
||(x_pointer == 25 && y_pointer == 100)
||(x_pointer == 26 && y_pointer == 100)
||(x_pointer == 27 && y_pointer == 100)
||(x_pointer == 28 && y_pointer == 100)
||(x_pointer == 29 && y_pointer == 100)
||(x_pointer == 30 && y_pointer == 100)
||(x_pointer == 31 && y_pointer == 100)
||(x_pointer == 32 && y_pointer == 100)
||(x_pointer == 33 && y_pointer == 100)
||(x_pointer == 34 && y_pointer == 100)
||(x_pointer == 35 && y_pointer == 100)
||(x_pointer == 36 && y_pointer == 100)
||(x_pointer == 37 && y_pointer == 100)
||(x_pointer == 38 && y_pointer == 100)
||(x_pointer == 39 && y_pointer == 100)
||(x_pointer == 40 && y_pointer == 100)
||(x_pointer == 41 && y_pointer == 100)
||(x_pointer == 42 && y_pointer == 100)
||(x_pointer == 43 && y_pointer == 100)
||(x_pointer == 122 && y_pointer == 100)
||(x_pointer == 123 && y_pointer == 100)
||(x_pointer == 124 && y_pointer == 100)
||(x_pointer == 125 && y_pointer == 100)
||(x_pointer == 126 && y_pointer == 100)
||(x_pointer == 127 && y_pointer == 100)
||(x_pointer == 128 && y_pointer == 100)
||(x_pointer == 129 && y_pointer == 100)
||(x_pointer == 130 && y_pointer == 100)
||(x_pointer == 131 && y_pointer == 100)
||(x_pointer == 132 && y_pointer == 100)
||(x_pointer == 133 && y_pointer == 100)
||(x_pointer == 134 && y_pointer == 100)
||(x_pointer == 135 && y_pointer == 100)
||(x_pointer == 136 && y_pointer == 100)
||(x_pointer == 137 && y_pointer == 100)
||(x_pointer == 138 && y_pointer == 100)
||(x_pointer == 139 && y_pointer == 100)
||(x_pointer == 140 && y_pointer == 100)
||(x_pointer == 141 && y_pointer == 100)
||(x_pointer == 142 && y_pointer == 100)
||(x_pointer == 23 && y_pointer == 101)
||(x_pointer == 24 && y_pointer == 101)
||(x_pointer == 25 && y_pointer == 101)
||(x_pointer == 26 && y_pointer == 101)
||(x_pointer == 27 && y_pointer == 101)
||(x_pointer == 28 && y_pointer == 101)
||(x_pointer == 29 && y_pointer == 101)
||(x_pointer == 30 && y_pointer == 101)
||(x_pointer == 31 && y_pointer == 101)
||(x_pointer == 32 && y_pointer == 101)
||(x_pointer == 33 && y_pointer == 101)
||(x_pointer == 34 && y_pointer == 101)
||(x_pointer == 35 && y_pointer == 101)
||(x_pointer == 36 && y_pointer == 101)
||(x_pointer == 37 && y_pointer == 101)
||(x_pointer == 38 && y_pointer == 101)
||(x_pointer == 39 && y_pointer == 101)
||(x_pointer == 40 && y_pointer == 101)
||(x_pointer == 41 && y_pointer == 101)
||(x_pointer == 42 && y_pointer == 101)
||(x_pointer == 43 && y_pointer == 101));


	wire barrier_pixel_4 = current_level == 4 && ((x_pointer == 32 && y_pointer == 5)
||(x_pointer == 33 && y_pointer == 5)
||(x_pointer == 34 && y_pointer == 5)
||(x_pointer == 35 && y_pointer == 5)
||(x_pointer == 36 && y_pointer == 5)
||(x_pointer == 37 && y_pointer == 5)
||(x_pointer == 38 && y_pointer == 5)
||(x_pointer == 39 && y_pointer == 5)
||(x_pointer == 40 && y_pointer == 5)
||(x_pointer == 32 && y_pointer == 6)
||(x_pointer == 33 && y_pointer == 6)
||(x_pointer == 34 && y_pointer == 6)
||(x_pointer == 35 && y_pointer == 6)
||(x_pointer == 36 && y_pointer == 6)
||(x_pointer == 37 && y_pointer == 6)
||(x_pointer == 38 && y_pointer == 6)
||(x_pointer == 39 && y_pointer == 6)
||(x_pointer == 40 && y_pointer == 6)
||(x_pointer == 32 && y_pointer == 7)
||(x_pointer == 33 && y_pointer == 7)
||(x_pointer == 34 && y_pointer == 7)
||(x_pointer == 35 && y_pointer == 7)
||(x_pointer == 36 && y_pointer == 7)
||(x_pointer == 37 && y_pointer == 7)
||(x_pointer == 38 && y_pointer == 7)
||(x_pointer == 39 && y_pointer == 7)
||(x_pointer == 40 && y_pointer == 7)
||(x_pointer == 32 && y_pointer == 8)
||(x_pointer == 33 && y_pointer == 8)
||(x_pointer == 34 && y_pointer == 8)
||(x_pointer == 35 && y_pointer == 8)
||(x_pointer == 36 && y_pointer == 8)
||(x_pointer == 37 && y_pointer == 8)
||(x_pointer == 38 && y_pointer == 8)
||(x_pointer == 39 && y_pointer == 8)
||(x_pointer == 40 && y_pointer == 8)
||(x_pointer == 32 && y_pointer == 9)
||(x_pointer == 33 && y_pointer == 9)
||(x_pointer == 34 && y_pointer == 9)
||(x_pointer == 35 && y_pointer == 9)
||(x_pointer == 36 && y_pointer == 9)
||(x_pointer == 37 && y_pointer == 9)
||(x_pointer == 38 && y_pointer == 9)
||(x_pointer == 39 && y_pointer == 9)
||(x_pointer == 40 && y_pointer == 9)
||(x_pointer == 32 && y_pointer == 10)
||(x_pointer == 33 && y_pointer == 10)
||(x_pointer == 34 && y_pointer == 10)
||(x_pointer == 35 && y_pointer == 10)
||(x_pointer == 36 && y_pointer == 10)
||(x_pointer == 37 && y_pointer == 10)
||(x_pointer == 38 && y_pointer == 10)
||(x_pointer == 39 && y_pointer == 10)
||(x_pointer == 40 && y_pointer == 10)
||(x_pointer == 32 && y_pointer == 11)
||(x_pointer == 33 && y_pointer == 11)
||(x_pointer == 34 && y_pointer == 11)
||(x_pointer == 35 && y_pointer == 11)
||(x_pointer == 36 && y_pointer == 11)
||(x_pointer == 37 && y_pointer == 11)
||(x_pointer == 38 && y_pointer == 11)
||(x_pointer == 39 && y_pointer == 11)
||(x_pointer == 40 && y_pointer == 11)
||(x_pointer == 32 && y_pointer == 12)
||(x_pointer == 33 && y_pointer == 12)
||(x_pointer == 34 && y_pointer == 12)
||(x_pointer == 35 && y_pointer == 12)
||(x_pointer == 36 && y_pointer == 12)
||(x_pointer == 37 && y_pointer == 12)
||(x_pointer == 38 && y_pointer == 12)
||(x_pointer == 39 && y_pointer == 12)
||(x_pointer == 40 && y_pointer == 12)
||(x_pointer == 32 && y_pointer == 13)
||(x_pointer == 33 && y_pointer == 13)
||(x_pointer == 34 && y_pointer == 13)
||(x_pointer == 35 && y_pointer == 13)
||(x_pointer == 36 && y_pointer == 13)
||(x_pointer == 37 && y_pointer == 13)
||(x_pointer == 38 && y_pointer == 13)
||(x_pointer == 39 && y_pointer == 13)
||(x_pointer == 40 && y_pointer == 13)
||(x_pointer == 32 && y_pointer == 14)
||(x_pointer == 33 && y_pointer == 14)
||(x_pointer == 34 && y_pointer == 14)
||(x_pointer == 35 && y_pointer == 14)
||(x_pointer == 36 && y_pointer == 14)
||(x_pointer == 37 && y_pointer == 14)
||(x_pointer == 38 && y_pointer == 14)
||(x_pointer == 39 && y_pointer == 14)
||(x_pointer == 40 && y_pointer == 14)
||(x_pointer == 32 && y_pointer == 15)
||(x_pointer == 33 && y_pointer == 15)
||(x_pointer == 34 && y_pointer == 15)
||(x_pointer == 35 && y_pointer == 15)
||(x_pointer == 36 && y_pointer == 15)
||(x_pointer == 37 && y_pointer == 15)
||(x_pointer == 38 && y_pointer == 15)
||(x_pointer == 39 && y_pointer == 15)
||(x_pointer == 40 && y_pointer == 15)
||(x_pointer == 32 && y_pointer == 16)
||(x_pointer == 33 && y_pointer == 16)
||(x_pointer == 34 && y_pointer == 16)
||(x_pointer == 35 && y_pointer == 16)
||(x_pointer == 36 && y_pointer == 16)
||(x_pointer == 37 && y_pointer == 16)
||(x_pointer == 38 && y_pointer == 16)
||(x_pointer == 39 && y_pointer == 16)
||(x_pointer == 40 && y_pointer == 16)
||(x_pointer == 32 && y_pointer == 17)
||(x_pointer == 33 && y_pointer == 17)
||(x_pointer == 34 && y_pointer == 17)
||(x_pointer == 35 && y_pointer == 17)
||(x_pointer == 36 && y_pointer == 17)
||(x_pointer == 37 && y_pointer == 17)
||(x_pointer == 38 && y_pointer == 17)
||(x_pointer == 39 && y_pointer == 17)
||(x_pointer == 40 && y_pointer == 17)
||(x_pointer == 32 && y_pointer == 18)
||(x_pointer == 33 && y_pointer == 18)
||(x_pointer == 34 && y_pointer == 18)
||(x_pointer == 35 && y_pointer == 18)
||(x_pointer == 36 && y_pointer == 18)
||(x_pointer == 37 && y_pointer == 18)
||(x_pointer == 38 && y_pointer == 18)
||(x_pointer == 39 && y_pointer == 18)
||(x_pointer == 40 && y_pointer == 18)
||(x_pointer == 32 && y_pointer == 19)
||(x_pointer == 33 && y_pointer == 19)
||(x_pointer == 34 && y_pointer == 19)
||(x_pointer == 35 && y_pointer == 19)
||(x_pointer == 36 && y_pointer == 19)
||(x_pointer == 37 && y_pointer == 19)
||(x_pointer == 38 && y_pointer == 19)
||(x_pointer == 39 && y_pointer == 19)
||(x_pointer == 40 && y_pointer == 19)
||(x_pointer == 32 && y_pointer == 20)
||(x_pointer == 33 && y_pointer == 20)
||(x_pointer == 34 && y_pointer == 20)
||(x_pointer == 35 && y_pointer == 20)
||(x_pointer == 36 && y_pointer == 20)
||(x_pointer == 37 && y_pointer == 20)
||(x_pointer == 38 && y_pointer == 20)
||(x_pointer == 39 && y_pointer == 20)
||(x_pointer == 40 && y_pointer == 20)
||(x_pointer == 32 && y_pointer == 21)
||(x_pointer == 33 && y_pointer == 21)
||(x_pointer == 34 && y_pointer == 21)
||(x_pointer == 35 && y_pointer == 21)
||(x_pointer == 36 && y_pointer == 21)
||(x_pointer == 37 && y_pointer == 21)
||(x_pointer == 38 && y_pointer == 21)
||(x_pointer == 39 && y_pointer == 21)
||(x_pointer == 40 && y_pointer == 21)
||(x_pointer == 32 && y_pointer == 22)
||(x_pointer == 33 && y_pointer == 22)
||(x_pointer == 34 && y_pointer == 22)
||(x_pointer == 35 && y_pointer == 22)
||(x_pointer == 36 && y_pointer == 22)
||(x_pointer == 37 && y_pointer == 22)
||(x_pointer == 38 && y_pointer == 22)
||(x_pointer == 39 && y_pointer == 22)
||(x_pointer == 40 && y_pointer == 22)
||(x_pointer == 32 && y_pointer == 23)
||(x_pointer == 33 && y_pointer == 23)
||(x_pointer == 34 && y_pointer == 23)
||(x_pointer == 35 && y_pointer == 23)
||(x_pointer == 36 && y_pointer == 23)
||(x_pointer == 37 && y_pointer == 23)
||(x_pointer == 38 && y_pointer == 23)
||(x_pointer == 39 && y_pointer == 23)
||(x_pointer == 40 && y_pointer == 23)
||(x_pointer == 32 && y_pointer == 24)
||(x_pointer == 33 && y_pointer == 24)
||(x_pointer == 34 && y_pointer == 24)
||(x_pointer == 35 && y_pointer == 24)
||(x_pointer == 36 && y_pointer == 24)
||(x_pointer == 37 && y_pointer == 24)
||(x_pointer == 38 && y_pointer == 24)
||(x_pointer == 39 && y_pointer == 24)
||(x_pointer == 40 && y_pointer == 24)
||(x_pointer == 32 && y_pointer == 25)
||(x_pointer == 33 && y_pointer == 25)
||(x_pointer == 34 && y_pointer == 25)
||(x_pointer == 35 && y_pointer == 25)
||(x_pointer == 36 && y_pointer == 25)
||(x_pointer == 37 && y_pointer == 25)
||(x_pointer == 38 && y_pointer == 25)
||(x_pointer == 39 && y_pointer == 25)
||(x_pointer == 40 && y_pointer == 25)
||(x_pointer == 32 && y_pointer == 26)
||(x_pointer == 33 && y_pointer == 26)
||(x_pointer == 34 && y_pointer == 26)
||(x_pointer == 35 && y_pointer == 26)
||(x_pointer == 36 && y_pointer == 26)
||(x_pointer == 37 && y_pointer == 26)
||(x_pointer == 38 && y_pointer == 26)
||(x_pointer == 39 && y_pointer == 26)
||(x_pointer == 40 && y_pointer == 26)
||(x_pointer == 32 && y_pointer == 27)
||(x_pointer == 33 && y_pointer == 27)
||(x_pointer == 34 && y_pointer == 27)
||(x_pointer == 35 && y_pointer == 27)
||(x_pointer == 36 && y_pointer == 27)
||(x_pointer == 37 && y_pointer == 27)
||(x_pointer == 38 && y_pointer == 27)
||(x_pointer == 39 && y_pointer == 27)
||(x_pointer == 40 && y_pointer == 27)
||(x_pointer == 32 && y_pointer == 28)
||(x_pointer == 33 && y_pointer == 28)
||(x_pointer == 34 && y_pointer == 28)
||(x_pointer == 35 && y_pointer == 28)
||(x_pointer == 36 && y_pointer == 28)
||(x_pointer == 37 && y_pointer == 28)
||(x_pointer == 38 && y_pointer == 28)
||(x_pointer == 39 && y_pointer == 28)
||(x_pointer == 40 && y_pointer == 28)
||(x_pointer == 32 && y_pointer == 29)
||(x_pointer == 33 && y_pointer == 29)
||(x_pointer == 34 && y_pointer == 29)
||(x_pointer == 35 && y_pointer == 29)
||(x_pointer == 36 && y_pointer == 29)
||(x_pointer == 37 && y_pointer == 29)
||(x_pointer == 38 && y_pointer == 29)
||(x_pointer == 39 && y_pointer == 29)
||(x_pointer == 40 && y_pointer == 29)
||(x_pointer == 32 && y_pointer == 30)
||(x_pointer == 33 && y_pointer == 30)
||(x_pointer == 34 && y_pointer == 30)
||(x_pointer == 35 && y_pointer == 30)
||(x_pointer == 36 && y_pointer == 30)
||(x_pointer == 37 && y_pointer == 30)
||(x_pointer == 38 && y_pointer == 30)
||(x_pointer == 39 && y_pointer == 30)
||(x_pointer == 40 && y_pointer == 30)
||(x_pointer == 32 && y_pointer == 31)
||(x_pointer == 33 && y_pointer == 31)
||(x_pointer == 34 && y_pointer == 31)
||(x_pointer == 35 && y_pointer == 31)
||(x_pointer == 36 && y_pointer == 31)
||(x_pointer == 37 && y_pointer == 31)
||(x_pointer == 38 && y_pointer == 31)
||(x_pointer == 39 && y_pointer == 31)
||(x_pointer == 40 && y_pointer == 31)
||(x_pointer == 32 && y_pointer == 32)
||(x_pointer == 33 && y_pointer == 32)
||(x_pointer == 34 && y_pointer == 32)
||(x_pointer == 35 && y_pointer == 32)
||(x_pointer == 36 && y_pointer == 32)
||(x_pointer == 37 && y_pointer == 32)
||(x_pointer == 38 && y_pointer == 32)
||(x_pointer == 39 && y_pointer == 32)
||(x_pointer == 40 && y_pointer == 32)
||(x_pointer == 32 && y_pointer == 33)
||(x_pointer == 33 && y_pointer == 33)
||(x_pointer == 34 && y_pointer == 33)
||(x_pointer == 35 && y_pointer == 33)
||(x_pointer == 36 && y_pointer == 33)
||(x_pointer == 37 && y_pointer == 33)
||(x_pointer == 38 && y_pointer == 33)
||(x_pointer == 39 && y_pointer == 33)
||(x_pointer == 40 && y_pointer == 33)
||(x_pointer == 32 && y_pointer == 34)
||(x_pointer == 33 && y_pointer == 34)
||(x_pointer == 34 && y_pointer == 34)
||(x_pointer == 35 && y_pointer == 34)
||(x_pointer == 36 && y_pointer == 34)
||(x_pointer == 37 && y_pointer == 34)
||(x_pointer == 38 && y_pointer == 34)
||(x_pointer == 39 && y_pointer == 34)
||(x_pointer == 40 && y_pointer == 34)
||(x_pointer == 32 && y_pointer == 35)
||(x_pointer == 33 && y_pointer == 35)
||(x_pointer == 34 && y_pointer == 35)
||(x_pointer == 35 && y_pointer == 35)
||(x_pointer == 36 && y_pointer == 35)
||(x_pointer == 37 && y_pointer == 35)
||(x_pointer == 38 && y_pointer == 35)
||(x_pointer == 39 && y_pointer == 35)
||(x_pointer == 40 && y_pointer == 35)
||(x_pointer == 32 && y_pointer == 36)
||(x_pointer == 33 && y_pointer == 36)
||(x_pointer == 34 && y_pointer == 36)
||(x_pointer == 35 && y_pointer == 36)
||(x_pointer == 36 && y_pointer == 36)
||(x_pointer == 37 && y_pointer == 36)
||(x_pointer == 38 && y_pointer == 36)
||(x_pointer == 39 && y_pointer == 36)
||(x_pointer == 40 && y_pointer == 36)
||(x_pointer == 32 && y_pointer == 37)
||(x_pointer == 33 && y_pointer == 37)
||(x_pointer == 34 && y_pointer == 37)
||(x_pointer == 35 && y_pointer == 37)
||(x_pointer == 36 && y_pointer == 37)
||(x_pointer == 37 && y_pointer == 37)
||(x_pointer == 38 && y_pointer == 37)
||(x_pointer == 39 && y_pointer == 37)
||(x_pointer == 40 && y_pointer == 37)
||(x_pointer == 32 && y_pointer == 38)
||(x_pointer == 33 && y_pointer == 38)
||(x_pointer == 34 && y_pointer == 38)
||(x_pointer == 35 && y_pointer == 38)
||(x_pointer == 36 && y_pointer == 38)
||(x_pointer == 37 && y_pointer == 38)
||(x_pointer == 38 && y_pointer == 38)
||(x_pointer == 39 && y_pointer == 38)
||(x_pointer == 40 && y_pointer == 38)
||(x_pointer == 71 && y_pointer == 38)
||(x_pointer == 72 && y_pointer == 38)
||(x_pointer == 73 && y_pointer == 38)
||(x_pointer == 74 && y_pointer == 38)
||(x_pointer == 75 && y_pointer == 38)
||(x_pointer == 76 && y_pointer == 38)
||(x_pointer == 77 && y_pointer == 38)
||(x_pointer == 78 && y_pointer == 38)
||(x_pointer == 79 && y_pointer == 38)
||(x_pointer == 80 && y_pointer == 38)
||(x_pointer == 81 && y_pointer == 38)
||(x_pointer == 82 && y_pointer == 38)
||(x_pointer == 83 && y_pointer == 38)
||(x_pointer == 84 && y_pointer == 38)
||(x_pointer == 85 && y_pointer == 38)
||(x_pointer == 86 && y_pointer == 38)
||(x_pointer == 87 && y_pointer == 38)
||(x_pointer == 88 && y_pointer == 38)
||(x_pointer == 89 && y_pointer == 38)
||(x_pointer == 90 && y_pointer == 38)
||(x_pointer == 91 && y_pointer == 38)
||(x_pointer == 92 && y_pointer == 38)
||(x_pointer == 93 && y_pointer == 38)
||(x_pointer == 94 && y_pointer == 38)
||(x_pointer == 95 && y_pointer == 38)
||(x_pointer == 96 && y_pointer == 38)
||(x_pointer == 97 && y_pointer == 38)
||(x_pointer == 98 && y_pointer == 38)
||(x_pointer == 99 && y_pointer == 38)
||(x_pointer == 100 && y_pointer == 38)
||(x_pointer == 101 && y_pointer == 38)
||(x_pointer == 102 && y_pointer == 38)
||(x_pointer == 103 && y_pointer == 38)
||(x_pointer == 104 && y_pointer == 38)
||(x_pointer == 105 && y_pointer == 38)
||(x_pointer == 106 && y_pointer == 38)
||(x_pointer == 107 && y_pointer == 38)
||(x_pointer == 108 && y_pointer == 38)
||(x_pointer == 109 && y_pointer == 38)
||(x_pointer == 110 && y_pointer == 38)
||(x_pointer == 111 && y_pointer == 38)
||(x_pointer == 112 && y_pointer == 38)
||(x_pointer == 113 && y_pointer == 38)
||(x_pointer == 114 && y_pointer == 38)
||(x_pointer == 115 && y_pointer == 38)
||(x_pointer == 116 && y_pointer == 38)
||(x_pointer == 117 && y_pointer == 38)
||(x_pointer == 118 && y_pointer == 38)
||(x_pointer == 119 && y_pointer == 38)
||(x_pointer == 120 && y_pointer == 38)
||(x_pointer == 121 && y_pointer == 38)
||(x_pointer == 122 && y_pointer == 38)
||(x_pointer == 123 && y_pointer == 38)
||(x_pointer == 124 && y_pointer == 38)
||(x_pointer == 125 && y_pointer == 38)
||(x_pointer == 126 && y_pointer == 38)
||(x_pointer == 127 && y_pointer == 38)
||(x_pointer == 128 && y_pointer == 38)
||(x_pointer == 129 && y_pointer == 38)
||(x_pointer == 130 && y_pointer == 38)
||(x_pointer == 131 && y_pointer == 38)
||(x_pointer == 132 && y_pointer == 38)
||(x_pointer == 133 && y_pointer == 38)
||(x_pointer == 134 && y_pointer == 38)
||(x_pointer == 135 && y_pointer == 38)
||(x_pointer == 136 && y_pointer == 38)
||(x_pointer == 137 && y_pointer == 38)
||(x_pointer == 138 && y_pointer == 38)
||(x_pointer == 139 && y_pointer == 38)
||(x_pointer == 140 && y_pointer == 38)
||(x_pointer == 141 && y_pointer == 38)
||(x_pointer == 142 && y_pointer == 38)
||(x_pointer == 143 && y_pointer == 38)
||(x_pointer == 144 && y_pointer == 38)
||(x_pointer == 145 && y_pointer == 38)
||(x_pointer == 146 && y_pointer == 38)
||(x_pointer == 147 && y_pointer == 38)
||(x_pointer == 148 && y_pointer == 38)
||(x_pointer == 149 && y_pointer == 38)
||(x_pointer == 150 && y_pointer == 38)
||(x_pointer == 151 && y_pointer == 38)
||(x_pointer == 152 && y_pointer == 38)
||(x_pointer == 153 && y_pointer == 38)
||(x_pointer == 154 && y_pointer == 38)
||(x_pointer == 32 && y_pointer == 39)
||(x_pointer == 33 && y_pointer == 39)
||(x_pointer == 34 && y_pointer == 39)
||(x_pointer == 35 && y_pointer == 39)
||(x_pointer == 36 && y_pointer == 39)
||(x_pointer == 37 && y_pointer == 39)
||(x_pointer == 38 && y_pointer == 39)
||(x_pointer == 39 && y_pointer == 39)
||(x_pointer == 40 && y_pointer == 39)
||(x_pointer == 71 && y_pointer == 39)
||(x_pointer == 72 && y_pointer == 39)
||(x_pointer == 73 && y_pointer == 39)
||(x_pointer == 74 && y_pointer == 39)
||(x_pointer == 75 && y_pointer == 39)
||(x_pointer == 76 && y_pointer == 39)
||(x_pointer == 77 && y_pointer == 39)
||(x_pointer == 78 && y_pointer == 39)
||(x_pointer == 79 && y_pointer == 39)
||(x_pointer == 80 && y_pointer == 39)
||(x_pointer == 81 && y_pointer == 39)
||(x_pointer == 82 && y_pointer == 39)
||(x_pointer == 83 && y_pointer == 39)
||(x_pointer == 84 && y_pointer == 39)
||(x_pointer == 85 && y_pointer == 39)
||(x_pointer == 86 && y_pointer == 39)
||(x_pointer == 87 && y_pointer == 39)
||(x_pointer == 88 && y_pointer == 39)
||(x_pointer == 89 && y_pointer == 39)
||(x_pointer == 90 && y_pointer == 39)
||(x_pointer == 91 && y_pointer == 39)
||(x_pointer == 92 && y_pointer == 39)
||(x_pointer == 93 && y_pointer == 39)
||(x_pointer == 94 && y_pointer == 39)
||(x_pointer == 95 && y_pointer == 39)
||(x_pointer == 96 && y_pointer == 39)
||(x_pointer == 97 && y_pointer == 39)
||(x_pointer == 98 && y_pointer == 39)
||(x_pointer == 99 && y_pointer == 39)
||(x_pointer == 100 && y_pointer == 39)
||(x_pointer == 101 && y_pointer == 39)
||(x_pointer == 102 && y_pointer == 39)
||(x_pointer == 103 && y_pointer == 39)
||(x_pointer == 104 && y_pointer == 39)
||(x_pointer == 105 && y_pointer == 39)
||(x_pointer == 106 && y_pointer == 39)
||(x_pointer == 107 && y_pointer == 39)
||(x_pointer == 108 && y_pointer == 39)
||(x_pointer == 109 && y_pointer == 39)
||(x_pointer == 110 && y_pointer == 39)
||(x_pointer == 111 && y_pointer == 39)
||(x_pointer == 112 && y_pointer == 39)
||(x_pointer == 113 && y_pointer == 39)
||(x_pointer == 114 && y_pointer == 39)
||(x_pointer == 115 && y_pointer == 39)
||(x_pointer == 116 && y_pointer == 39)
||(x_pointer == 117 && y_pointer == 39)
||(x_pointer == 118 && y_pointer == 39)
||(x_pointer == 119 && y_pointer == 39)
||(x_pointer == 120 && y_pointer == 39)
||(x_pointer == 121 && y_pointer == 39)
||(x_pointer == 122 && y_pointer == 39)
||(x_pointer == 123 && y_pointer == 39)
||(x_pointer == 124 && y_pointer == 39)
||(x_pointer == 125 && y_pointer == 39)
||(x_pointer == 126 && y_pointer == 39)
||(x_pointer == 127 && y_pointer == 39)
||(x_pointer == 128 && y_pointer == 39)
||(x_pointer == 129 && y_pointer == 39)
||(x_pointer == 130 && y_pointer == 39)
||(x_pointer == 131 && y_pointer == 39)
||(x_pointer == 132 && y_pointer == 39)
||(x_pointer == 133 && y_pointer == 39)
||(x_pointer == 134 && y_pointer == 39)
||(x_pointer == 135 && y_pointer == 39)
||(x_pointer == 136 && y_pointer == 39)
||(x_pointer == 137 && y_pointer == 39)
||(x_pointer == 138 && y_pointer == 39)
||(x_pointer == 139 && y_pointer == 39)
||(x_pointer == 140 && y_pointer == 39)
||(x_pointer == 141 && y_pointer == 39)
||(x_pointer == 142 && y_pointer == 39)
||(x_pointer == 143 && y_pointer == 39)
||(x_pointer == 144 && y_pointer == 39)
||(x_pointer == 145 && y_pointer == 39)
||(x_pointer == 146 && y_pointer == 39)
||(x_pointer == 147 && y_pointer == 39)
||(x_pointer == 148 && y_pointer == 39)
||(x_pointer == 149 && y_pointer == 39)
||(x_pointer == 150 && y_pointer == 39)
||(x_pointer == 151 && y_pointer == 39)
||(x_pointer == 152 && y_pointer == 39)
||(x_pointer == 153 && y_pointer == 39)
||(x_pointer == 154 && y_pointer == 39)
||(x_pointer == 32 && y_pointer == 40)
||(x_pointer == 33 && y_pointer == 40)
||(x_pointer == 34 && y_pointer == 40)
||(x_pointer == 35 && y_pointer == 40)
||(x_pointer == 36 && y_pointer == 40)
||(x_pointer == 37 && y_pointer == 40)
||(x_pointer == 38 && y_pointer == 40)
||(x_pointer == 39 && y_pointer == 40)
||(x_pointer == 40 && y_pointer == 40)
||(x_pointer == 71 && y_pointer == 40)
||(x_pointer == 72 && y_pointer == 40)
||(x_pointer == 73 && y_pointer == 40)
||(x_pointer == 74 && y_pointer == 40)
||(x_pointer == 75 && y_pointer == 40)
||(x_pointer == 76 && y_pointer == 40)
||(x_pointer == 77 && y_pointer == 40)
||(x_pointer == 78 && y_pointer == 40)
||(x_pointer == 79 && y_pointer == 40)
||(x_pointer == 80 && y_pointer == 40)
||(x_pointer == 81 && y_pointer == 40)
||(x_pointer == 82 && y_pointer == 40)
||(x_pointer == 83 && y_pointer == 40)
||(x_pointer == 84 && y_pointer == 40)
||(x_pointer == 85 && y_pointer == 40)
||(x_pointer == 86 && y_pointer == 40)
||(x_pointer == 87 && y_pointer == 40)
||(x_pointer == 88 && y_pointer == 40)
||(x_pointer == 89 && y_pointer == 40)
||(x_pointer == 90 && y_pointer == 40)
||(x_pointer == 91 && y_pointer == 40)
||(x_pointer == 92 && y_pointer == 40)
||(x_pointer == 93 && y_pointer == 40)
||(x_pointer == 94 && y_pointer == 40)
||(x_pointer == 95 && y_pointer == 40)
||(x_pointer == 96 && y_pointer == 40)
||(x_pointer == 97 && y_pointer == 40)
||(x_pointer == 98 && y_pointer == 40)
||(x_pointer == 99 && y_pointer == 40)
||(x_pointer == 100 && y_pointer == 40)
||(x_pointer == 101 && y_pointer == 40)
||(x_pointer == 102 && y_pointer == 40)
||(x_pointer == 103 && y_pointer == 40)
||(x_pointer == 104 && y_pointer == 40)
||(x_pointer == 105 && y_pointer == 40)
||(x_pointer == 106 && y_pointer == 40)
||(x_pointer == 107 && y_pointer == 40)
||(x_pointer == 108 && y_pointer == 40)
||(x_pointer == 109 && y_pointer == 40)
||(x_pointer == 110 && y_pointer == 40)
||(x_pointer == 111 && y_pointer == 40)
||(x_pointer == 112 && y_pointer == 40)
||(x_pointer == 113 && y_pointer == 40)
||(x_pointer == 114 && y_pointer == 40)
||(x_pointer == 115 && y_pointer == 40)
||(x_pointer == 116 && y_pointer == 40)
||(x_pointer == 117 && y_pointer == 40)
||(x_pointer == 118 && y_pointer == 40)
||(x_pointer == 119 && y_pointer == 40)
||(x_pointer == 120 && y_pointer == 40)
||(x_pointer == 121 && y_pointer == 40)
||(x_pointer == 122 && y_pointer == 40)
||(x_pointer == 123 && y_pointer == 40)
||(x_pointer == 124 && y_pointer == 40)
||(x_pointer == 125 && y_pointer == 40)
||(x_pointer == 126 && y_pointer == 40)
||(x_pointer == 127 && y_pointer == 40)
||(x_pointer == 128 && y_pointer == 40)
||(x_pointer == 129 && y_pointer == 40)
||(x_pointer == 130 && y_pointer == 40)
||(x_pointer == 131 && y_pointer == 40)
||(x_pointer == 132 && y_pointer == 40)
||(x_pointer == 133 && y_pointer == 40)
||(x_pointer == 134 && y_pointer == 40)
||(x_pointer == 135 && y_pointer == 40)
||(x_pointer == 136 && y_pointer == 40)
||(x_pointer == 137 && y_pointer == 40)
||(x_pointer == 138 && y_pointer == 40)
||(x_pointer == 139 && y_pointer == 40)
||(x_pointer == 140 && y_pointer == 40)
||(x_pointer == 141 && y_pointer == 40)
||(x_pointer == 142 && y_pointer == 40)
||(x_pointer == 143 && y_pointer == 40)
||(x_pointer == 144 && y_pointer == 40)
||(x_pointer == 145 && y_pointer == 40)
||(x_pointer == 146 && y_pointer == 40)
||(x_pointer == 147 && y_pointer == 40)
||(x_pointer == 148 && y_pointer == 40)
||(x_pointer == 149 && y_pointer == 40)
||(x_pointer == 150 && y_pointer == 40)
||(x_pointer == 151 && y_pointer == 40)
||(x_pointer == 152 && y_pointer == 40)
||(x_pointer == 153 && y_pointer == 40)
||(x_pointer == 154 && y_pointer == 40)
||(x_pointer == 32 && y_pointer == 41)
||(x_pointer == 33 && y_pointer == 41)
||(x_pointer == 34 && y_pointer == 41)
||(x_pointer == 35 && y_pointer == 41)
||(x_pointer == 36 && y_pointer == 41)
||(x_pointer == 37 && y_pointer == 41)
||(x_pointer == 38 && y_pointer == 41)
||(x_pointer == 39 && y_pointer == 41)
||(x_pointer == 40 && y_pointer == 41)
||(x_pointer == 71 && y_pointer == 41)
||(x_pointer == 72 && y_pointer == 41)
||(x_pointer == 73 && y_pointer == 41)
||(x_pointer == 74 && y_pointer == 41)
||(x_pointer == 75 && y_pointer == 41)
||(x_pointer == 76 && y_pointer == 41)
||(x_pointer == 77 && y_pointer == 41)
||(x_pointer == 78 && y_pointer == 41)
||(x_pointer == 79 && y_pointer == 41)
||(x_pointer == 80 && y_pointer == 41)
||(x_pointer == 81 && y_pointer == 41)
||(x_pointer == 82 && y_pointer == 41)
||(x_pointer == 83 && y_pointer == 41)
||(x_pointer == 84 && y_pointer == 41)
||(x_pointer == 85 && y_pointer == 41)
||(x_pointer == 86 && y_pointer == 41)
||(x_pointer == 87 && y_pointer == 41)
||(x_pointer == 88 && y_pointer == 41)
||(x_pointer == 89 && y_pointer == 41)
||(x_pointer == 90 && y_pointer == 41)
||(x_pointer == 91 && y_pointer == 41)
||(x_pointer == 92 && y_pointer == 41)
||(x_pointer == 93 && y_pointer == 41)
||(x_pointer == 94 && y_pointer == 41)
||(x_pointer == 95 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 99 && y_pointer == 41)
||(x_pointer == 100 && y_pointer == 41)
||(x_pointer == 101 && y_pointer == 41)
||(x_pointer == 102 && y_pointer == 41)
||(x_pointer == 103 && y_pointer == 41)
||(x_pointer == 104 && y_pointer == 41)
||(x_pointer == 105 && y_pointer == 41)
||(x_pointer == 106 && y_pointer == 41)
||(x_pointer == 107 && y_pointer == 41)
||(x_pointer == 108 && y_pointer == 41)
||(x_pointer == 109 && y_pointer == 41)
||(x_pointer == 110 && y_pointer == 41)
||(x_pointer == 111 && y_pointer == 41)
||(x_pointer == 112 && y_pointer == 41)
||(x_pointer == 113 && y_pointer == 41)
||(x_pointer == 114 && y_pointer == 41)
||(x_pointer == 115 && y_pointer == 41)
||(x_pointer == 116 && y_pointer == 41)
||(x_pointer == 117 && y_pointer == 41)
||(x_pointer == 118 && y_pointer == 41)
||(x_pointer == 119 && y_pointer == 41)
||(x_pointer == 120 && y_pointer == 41)
||(x_pointer == 121 && y_pointer == 41)
||(x_pointer == 122 && y_pointer == 41)
||(x_pointer == 123 && y_pointer == 41)
||(x_pointer == 124 && y_pointer == 41)
||(x_pointer == 125 && y_pointer == 41)
||(x_pointer == 126 && y_pointer == 41)
||(x_pointer == 127 && y_pointer == 41)
||(x_pointer == 128 && y_pointer == 41)
||(x_pointer == 129 && y_pointer == 41)
||(x_pointer == 130 && y_pointer == 41)
||(x_pointer == 131 && y_pointer == 41)
||(x_pointer == 132 && y_pointer == 41)
||(x_pointer == 133 && y_pointer == 41)
||(x_pointer == 134 && y_pointer == 41)
||(x_pointer == 135 && y_pointer == 41)
||(x_pointer == 136 && y_pointer == 41)
||(x_pointer == 137 && y_pointer == 41)
||(x_pointer == 138 && y_pointer == 41)
||(x_pointer == 139 && y_pointer == 41)
||(x_pointer == 140 && y_pointer == 41)
||(x_pointer == 141 && y_pointer == 41)
||(x_pointer == 142 && y_pointer == 41)
||(x_pointer == 143 && y_pointer == 41)
||(x_pointer == 144 && y_pointer == 41)
||(x_pointer == 145 && y_pointer == 41)
||(x_pointer == 146 && y_pointer == 41)
||(x_pointer == 147 && y_pointer == 41)
||(x_pointer == 148 && y_pointer == 41)
||(x_pointer == 149 && y_pointer == 41)
||(x_pointer == 150 && y_pointer == 41)
||(x_pointer == 151 && y_pointer == 41)
||(x_pointer == 152 && y_pointer == 41)
||(x_pointer == 153 && y_pointer == 41)
||(x_pointer == 154 && y_pointer == 41)
||(x_pointer == 32 && y_pointer == 42)
||(x_pointer == 33 && y_pointer == 42)
||(x_pointer == 34 && y_pointer == 42)
||(x_pointer == 35 && y_pointer == 42)
||(x_pointer == 36 && y_pointer == 42)
||(x_pointer == 37 && y_pointer == 42)
||(x_pointer == 38 && y_pointer == 42)
||(x_pointer == 39 && y_pointer == 42)
||(x_pointer == 40 && y_pointer == 42)
||(x_pointer == 71 && y_pointer == 42)
||(x_pointer == 72 && y_pointer == 42)
||(x_pointer == 73 && y_pointer == 42)
||(x_pointer == 74 && y_pointer == 42)
||(x_pointer == 75 && y_pointer == 42)
||(x_pointer == 76 && y_pointer == 42)
||(x_pointer == 77 && y_pointer == 42)
||(x_pointer == 78 && y_pointer == 42)
||(x_pointer == 79 && y_pointer == 42)
||(x_pointer == 80 && y_pointer == 42)
||(x_pointer == 81 && y_pointer == 42)
||(x_pointer == 82 && y_pointer == 42)
||(x_pointer == 83 && y_pointer == 42)
||(x_pointer == 84 && y_pointer == 42)
||(x_pointer == 85 && y_pointer == 42)
||(x_pointer == 86 && y_pointer == 42)
||(x_pointer == 87 && y_pointer == 42)
||(x_pointer == 88 && y_pointer == 42)
||(x_pointer == 89 && y_pointer == 42)
||(x_pointer == 90 && y_pointer == 42)
||(x_pointer == 91 && y_pointer == 42)
||(x_pointer == 92 && y_pointer == 42)
||(x_pointer == 93 && y_pointer == 42)
||(x_pointer == 94 && y_pointer == 42)
||(x_pointer == 95 && y_pointer == 42)
||(x_pointer == 96 && y_pointer == 42)
||(x_pointer == 97 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 99 && y_pointer == 42)
||(x_pointer == 100 && y_pointer == 42)
||(x_pointer == 101 && y_pointer == 42)
||(x_pointer == 102 && y_pointer == 42)
||(x_pointer == 103 && y_pointer == 42)
||(x_pointer == 104 && y_pointer == 42)
||(x_pointer == 105 && y_pointer == 42)
||(x_pointer == 106 && y_pointer == 42)
||(x_pointer == 107 && y_pointer == 42)
||(x_pointer == 108 && y_pointer == 42)
||(x_pointer == 109 && y_pointer == 42)
||(x_pointer == 110 && y_pointer == 42)
||(x_pointer == 111 && y_pointer == 42)
||(x_pointer == 112 && y_pointer == 42)
||(x_pointer == 113 && y_pointer == 42)
||(x_pointer == 114 && y_pointer == 42)
||(x_pointer == 115 && y_pointer == 42)
||(x_pointer == 116 && y_pointer == 42)
||(x_pointer == 117 && y_pointer == 42)
||(x_pointer == 118 && y_pointer == 42)
||(x_pointer == 119 && y_pointer == 42)
||(x_pointer == 120 && y_pointer == 42)
||(x_pointer == 121 && y_pointer == 42)
||(x_pointer == 122 && y_pointer == 42)
||(x_pointer == 123 && y_pointer == 42)
||(x_pointer == 124 && y_pointer == 42)
||(x_pointer == 125 && y_pointer == 42)
||(x_pointer == 126 && y_pointer == 42)
||(x_pointer == 127 && y_pointer == 42)
||(x_pointer == 128 && y_pointer == 42)
||(x_pointer == 129 && y_pointer == 42)
||(x_pointer == 130 && y_pointer == 42)
||(x_pointer == 131 && y_pointer == 42)
||(x_pointer == 132 && y_pointer == 42)
||(x_pointer == 133 && y_pointer == 42)
||(x_pointer == 134 && y_pointer == 42)
||(x_pointer == 135 && y_pointer == 42)
||(x_pointer == 136 && y_pointer == 42)
||(x_pointer == 137 && y_pointer == 42)
||(x_pointer == 138 && y_pointer == 42)
||(x_pointer == 139 && y_pointer == 42)
||(x_pointer == 140 && y_pointer == 42)
||(x_pointer == 141 && y_pointer == 42)
||(x_pointer == 142 && y_pointer == 42)
||(x_pointer == 143 && y_pointer == 42)
||(x_pointer == 144 && y_pointer == 42)
||(x_pointer == 145 && y_pointer == 42)
||(x_pointer == 146 && y_pointer == 42)
||(x_pointer == 147 && y_pointer == 42)
||(x_pointer == 148 && y_pointer == 42)
||(x_pointer == 149 && y_pointer == 42)
||(x_pointer == 150 && y_pointer == 42)
||(x_pointer == 151 && y_pointer == 42)
||(x_pointer == 152 && y_pointer == 42)
||(x_pointer == 153 && y_pointer == 42)
||(x_pointer == 154 && y_pointer == 42)
||(x_pointer == 32 && y_pointer == 43)
||(x_pointer == 33 && y_pointer == 43)
||(x_pointer == 34 && y_pointer == 43)
||(x_pointer == 35 && y_pointer == 43)
||(x_pointer == 36 && y_pointer == 43)
||(x_pointer == 37 && y_pointer == 43)
||(x_pointer == 38 && y_pointer == 43)
||(x_pointer == 39 && y_pointer == 43)
||(x_pointer == 40 && y_pointer == 43)
||(x_pointer == 71 && y_pointer == 43)
||(x_pointer == 72 && y_pointer == 43)
||(x_pointer == 73 && y_pointer == 43)
||(x_pointer == 74 && y_pointer == 43)
||(x_pointer == 75 && y_pointer == 43)
||(x_pointer == 76 && y_pointer == 43)
||(x_pointer == 77 && y_pointer == 43)
||(x_pointer == 78 && y_pointer == 43)
||(x_pointer == 79 && y_pointer == 43)
||(x_pointer == 80 && y_pointer == 43)
||(x_pointer == 81 && y_pointer == 43)
||(x_pointer == 82 && y_pointer == 43)
||(x_pointer == 83 && y_pointer == 43)
||(x_pointer == 84 && y_pointer == 43)
||(x_pointer == 85 && y_pointer == 43)
||(x_pointer == 86 && y_pointer == 43)
||(x_pointer == 87 && y_pointer == 43)
||(x_pointer == 88 && y_pointer == 43)
||(x_pointer == 89 && y_pointer == 43)
||(x_pointer == 90 && y_pointer == 43)
||(x_pointer == 91 && y_pointer == 43)
||(x_pointer == 92 && y_pointer == 43)
||(x_pointer == 93 && y_pointer == 43)
||(x_pointer == 94 && y_pointer == 43)
||(x_pointer == 95 && y_pointer == 43)
||(x_pointer == 96 && y_pointer == 43)
||(x_pointer == 97 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 99 && y_pointer == 43)
||(x_pointer == 100 && y_pointer == 43)
||(x_pointer == 101 && y_pointer == 43)
||(x_pointer == 102 && y_pointer == 43)
||(x_pointer == 103 && y_pointer == 43)
||(x_pointer == 104 && y_pointer == 43)
||(x_pointer == 105 && y_pointer == 43)
||(x_pointer == 106 && y_pointer == 43)
||(x_pointer == 107 && y_pointer == 43)
||(x_pointer == 108 && y_pointer == 43)
||(x_pointer == 109 && y_pointer == 43)
||(x_pointer == 110 && y_pointer == 43)
||(x_pointer == 111 && y_pointer == 43)
||(x_pointer == 112 && y_pointer == 43)
||(x_pointer == 113 && y_pointer == 43)
||(x_pointer == 114 && y_pointer == 43)
||(x_pointer == 115 && y_pointer == 43)
||(x_pointer == 116 && y_pointer == 43)
||(x_pointer == 117 && y_pointer == 43)
||(x_pointer == 118 && y_pointer == 43)
||(x_pointer == 119 && y_pointer == 43)
||(x_pointer == 120 && y_pointer == 43)
||(x_pointer == 121 && y_pointer == 43)
||(x_pointer == 122 && y_pointer == 43)
||(x_pointer == 123 && y_pointer == 43)
||(x_pointer == 124 && y_pointer == 43)
||(x_pointer == 125 && y_pointer == 43)
||(x_pointer == 126 && y_pointer == 43)
||(x_pointer == 127 && y_pointer == 43)
||(x_pointer == 128 && y_pointer == 43)
||(x_pointer == 129 && y_pointer == 43)
||(x_pointer == 130 && y_pointer == 43)
||(x_pointer == 131 && y_pointer == 43)
||(x_pointer == 132 && y_pointer == 43)
||(x_pointer == 133 && y_pointer == 43)
||(x_pointer == 134 && y_pointer == 43)
||(x_pointer == 135 && y_pointer == 43)
||(x_pointer == 136 && y_pointer == 43)
||(x_pointer == 137 && y_pointer == 43)
||(x_pointer == 138 && y_pointer == 43)
||(x_pointer == 139 && y_pointer == 43)
||(x_pointer == 140 && y_pointer == 43)
||(x_pointer == 141 && y_pointer == 43)
||(x_pointer == 142 && y_pointer == 43)
||(x_pointer == 143 && y_pointer == 43)
||(x_pointer == 144 && y_pointer == 43)
||(x_pointer == 145 && y_pointer == 43)
||(x_pointer == 146 && y_pointer == 43)
||(x_pointer == 147 && y_pointer == 43)
||(x_pointer == 148 && y_pointer == 43)
||(x_pointer == 149 && y_pointer == 43)
||(x_pointer == 150 && y_pointer == 43)
||(x_pointer == 151 && y_pointer == 43)
||(x_pointer == 152 && y_pointer == 43)
||(x_pointer == 153 && y_pointer == 43)
||(x_pointer == 154 && y_pointer == 43)
||(x_pointer == 32 && y_pointer == 44)
||(x_pointer == 33 && y_pointer == 44)
||(x_pointer == 34 && y_pointer == 44)
||(x_pointer == 35 && y_pointer == 44)
||(x_pointer == 36 && y_pointer == 44)
||(x_pointer == 37 && y_pointer == 44)
||(x_pointer == 38 && y_pointer == 44)
||(x_pointer == 39 && y_pointer == 44)
||(x_pointer == 40 && y_pointer == 44)
||(x_pointer == 71 && y_pointer == 44)
||(x_pointer == 72 && y_pointer == 44)
||(x_pointer == 73 && y_pointer == 44)
||(x_pointer == 74 && y_pointer == 44)
||(x_pointer == 75 && y_pointer == 44)
||(x_pointer == 76 && y_pointer == 44)
||(x_pointer == 77 && y_pointer == 44)
||(x_pointer == 78 && y_pointer == 44)
||(x_pointer == 79 && y_pointer == 44)
||(x_pointer == 80 && y_pointer == 44)
||(x_pointer == 81 && y_pointer == 44)
||(x_pointer == 82 && y_pointer == 44)
||(x_pointer == 83 && y_pointer == 44)
||(x_pointer == 84 && y_pointer == 44)
||(x_pointer == 85 && y_pointer == 44)
||(x_pointer == 86 && y_pointer == 44)
||(x_pointer == 87 && y_pointer == 44)
||(x_pointer == 88 && y_pointer == 44)
||(x_pointer == 89 && y_pointer == 44)
||(x_pointer == 90 && y_pointer == 44)
||(x_pointer == 91 && y_pointer == 44)
||(x_pointer == 92 && y_pointer == 44)
||(x_pointer == 93 && y_pointer == 44)
||(x_pointer == 94 && y_pointer == 44)
||(x_pointer == 95 && y_pointer == 44)
||(x_pointer == 96 && y_pointer == 44)
||(x_pointer == 97 && y_pointer == 44)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 99 && y_pointer == 44)
||(x_pointer == 100 && y_pointer == 44)
||(x_pointer == 101 && y_pointer == 44)
||(x_pointer == 102 && y_pointer == 44)
||(x_pointer == 103 && y_pointer == 44)
||(x_pointer == 104 && y_pointer == 44)
||(x_pointer == 105 && y_pointer == 44)
||(x_pointer == 106 && y_pointer == 44)
||(x_pointer == 107 && y_pointer == 44)
||(x_pointer == 108 && y_pointer == 44)
||(x_pointer == 109 && y_pointer == 44)
||(x_pointer == 110 && y_pointer == 44)
||(x_pointer == 111 && y_pointer == 44)
||(x_pointer == 112 && y_pointer == 44)
||(x_pointer == 113 && y_pointer == 44)
||(x_pointer == 114 && y_pointer == 44)
||(x_pointer == 115 && y_pointer == 44)
||(x_pointer == 116 && y_pointer == 44)
||(x_pointer == 117 && y_pointer == 44)
||(x_pointer == 118 && y_pointer == 44)
||(x_pointer == 119 && y_pointer == 44)
||(x_pointer == 120 && y_pointer == 44)
||(x_pointer == 121 && y_pointer == 44)
||(x_pointer == 122 && y_pointer == 44)
||(x_pointer == 123 && y_pointer == 44)
||(x_pointer == 124 && y_pointer == 44)
||(x_pointer == 125 && y_pointer == 44)
||(x_pointer == 126 && y_pointer == 44)
||(x_pointer == 127 && y_pointer == 44)
||(x_pointer == 128 && y_pointer == 44)
||(x_pointer == 129 && y_pointer == 44)
||(x_pointer == 130 && y_pointer == 44)
||(x_pointer == 131 && y_pointer == 44)
||(x_pointer == 132 && y_pointer == 44)
||(x_pointer == 133 && y_pointer == 44)
||(x_pointer == 134 && y_pointer == 44)
||(x_pointer == 135 && y_pointer == 44)
||(x_pointer == 136 && y_pointer == 44)
||(x_pointer == 137 && y_pointer == 44)
||(x_pointer == 138 && y_pointer == 44)
||(x_pointer == 139 && y_pointer == 44)
||(x_pointer == 140 && y_pointer == 44)
||(x_pointer == 141 && y_pointer == 44)
||(x_pointer == 142 && y_pointer == 44)
||(x_pointer == 143 && y_pointer == 44)
||(x_pointer == 144 && y_pointer == 44)
||(x_pointer == 145 && y_pointer == 44)
||(x_pointer == 146 && y_pointer == 44)
||(x_pointer == 147 && y_pointer == 44)
||(x_pointer == 148 && y_pointer == 44)
||(x_pointer == 149 && y_pointer == 44)
||(x_pointer == 150 && y_pointer == 44)
||(x_pointer == 151 && y_pointer == 44)
||(x_pointer == 152 && y_pointer == 44)
||(x_pointer == 153 && y_pointer == 44)
||(x_pointer == 154 && y_pointer == 44)
||(x_pointer == 32 && y_pointer == 45)
||(x_pointer == 33 && y_pointer == 45)
||(x_pointer == 34 && y_pointer == 45)
||(x_pointer == 35 && y_pointer == 45)
||(x_pointer == 36 && y_pointer == 45)
||(x_pointer == 37 && y_pointer == 45)
||(x_pointer == 38 && y_pointer == 45)
||(x_pointer == 39 && y_pointer == 45)
||(x_pointer == 40 && y_pointer == 45)
||(x_pointer == 71 && y_pointer == 45)
||(x_pointer == 72 && y_pointer == 45)
||(x_pointer == 73 && y_pointer == 45)
||(x_pointer == 74 && y_pointer == 45)
||(x_pointer == 75 && y_pointer == 45)
||(x_pointer == 76 && y_pointer == 45)
||(x_pointer == 77 && y_pointer == 45)
||(x_pointer == 78 && y_pointer == 45)
||(x_pointer == 79 && y_pointer == 45)
||(x_pointer == 80 && y_pointer == 45)
||(x_pointer == 81 && y_pointer == 45)
||(x_pointer == 82 && y_pointer == 45)
||(x_pointer == 83 && y_pointer == 45)
||(x_pointer == 84 && y_pointer == 45)
||(x_pointer == 85 && y_pointer == 45)
||(x_pointer == 86 && y_pointer == 45)
||(x_pointer == 87 && y_pointer == 45)
||(x_pointer == 88 && y_pointer == 45)
||(x_pointer == 89 && y_pointer == 45)
||(x_pointer == 90 && y_pointer == 45)
||(x_pointer == 91 && y_pointer == 45)
||(x_pointer == 92 && y_pointer == 45)
||(x_pointer == 93 && y_pointer == 45)
||(x_pointer == 94 && y_pointer == 45)
||(x_pointer == 95 && y_pointer == 45)
||(x_pointer == 96 && y_pointer == 45)
||(x_pointer == 97 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 99 && y_pointer == 45)
||(x_pointer == 100 && y_pointer == 45)
||(x_pointer == 101 && y_pointer == 45)
||(x_pointer == 102 && y_pointer == 45)
||(x_pointer == 103 && y_pointer == 45)
||(x_pointer == 104 && y_pointer == 45)
||(x_pointer == 105 && y_pointer == 45)
||(x_pointer == 106 && y_pointer == 45)
||(x_pointer == 107 && y_pointer == 45)
||(x_pointer == 108 && y_pointer == 45)
||(x_pointer == 109 && y_pointer == 45)
||(x_pointer == 110 && y_pointer == 45)
||(x_pointer == 111 && y_pointer == 45)
||(x_pointer == 112 && y_pointer == 45)
||(x_pointer == 113 && y_pointer == 45)
||(x_pointer == 114 && y_pointer == 45)
||(x_pointer == 115 && y_pointer == 45)
||(x_pointer == 116 && y_pointer == 45)
||(x_pointer == 117 && y_pointer == 45)
||(x_pointer == 118 && y_pointer == 45)
||(x_pointer == 119 && y_pointer == 45)
||(x_pointer == 120 && y_pointer == 45)
||(x_pointer == 121 && y_pointer == 45)
||(x_pointer == 122 && y_pointer == 45)
||(x_pointer == 123 && y_pointer == 45)
||(x_pointer == 124 && y_pointer == 45)
||(x_pointer == 125 && y_pointer == 45)
||(x_pointer == 126 && y_pointer == 45)
||(x_pointer == 127 && y_pointer == 45)
||(x_pointer == 128 && y_pointer == 45)
||(x_pointer == 129 && y_pointer == 45)
||(x_pointer == 130 && y_pointer == 45)
||(x_pointer == 131 && y_pointer == 45)
||(x_pointer == 132 && y_pointer == 45)
||(x_pointer == 133 && y_pointer == 45)
||(x_pointer == 134 && y_pointer == 45)
||(x_pointer == 135 && y_pointer == 45)
||(x_pointer == 136 && y_pointer == 45)
||(x_pointer == 137 && y_pointer == 45)
||(x_pointer == 138 && y_pointer == 45)
||(x_pointer == 139 && y_pointer == 45)
||(x_pointer == 140 && y_pointer == 45)
||(x_pointer == 141 && y_pointer == 45)
||(x_pointer == 142 && y_pointer == 45)
||(x_pointer == 143 && y_pointer == 45)
||(x_pointer == 144 && y_pointer == 45)
||(x_pointer == 145 && y_pointer == 45)
||(x_pointer == 146 && y_pointer == 45)
||(x_pointer == 147 && y_pointer == 45)
||(x_pointer == 148 && y_pointer == 45)
||(x_pointer == 149 && y_pointer == 45)
||(x_pointer == 150 && y_pointer == 45)
||(x_pointer == 151 && y_pointer == 45)
||(x_pointer == 152 && y_pointer == 45)
||(x_pointer == 153 && y_pointer == 45)
||(x_pointer == 154 && y_pointer == 45)
||(x_pointer == 32 && y_pointer == 46)
||(x_pointer == 33 && y_pointer == 46)
||(x_pointer == 34 && y_pointer == 46)
||(x_pointer == 35 && y_pointer == 46)
||(x_pointer == 36 && y_pointer == 46)
||(x_pointer == 37 && y_pointer == 46)
||(x_pointer == 38 && y_pointer == 46)
||(x_pointer == 39 && y_pointer == 46)
||(x_pointer == 40 && y_pointer == 46)
||(x_pointer == 71 && y_pointer == 46)
||(x_pointer == 72 && y_pointer == 46)
||(x_pointer == 73 && y_pointer == 46)
||(x_pointer == 74 && y_pointer == 46)
||(x_pointer == 75 && y_pointer == 46)
||(x_pointer == 76 && y_pointer == 46)
||(x_pointer == 77 && y_pointer == 46)
||(x_pointer == 78 && y_pointer == 46)
||(x_pointer == 79 && y_pointer == 46)
||(x_pointer == 80 && y_pointer == 46)
||(x_pointer == 81 && y_pointer == 46)
||(x_pointer == 82 && y_pointer == 46)
||(x_pointer == 83 && y_pointer == 46)
||(x_pointer == 84 && y_pointer == 46)
||(x_pointer == 85 && y_pointer == 46)
||(x_pointer == 86 && y_pointer == 46)
||(x_pointer == 87 && y_pointer == 46)
||(x_pointer == 88 && y_pointer == 46)
||(x_pointer == 89 && y_pointer == 46)
||(x_pointer == 90 && y_pointer == 46)
||(x_pointer == 91 && y_pointer == 46)
||(x_pointer == 92 && y_pointer == 46)
||(x_pointer == 93 && y_pointer == 46)
||(x_pointer == 94 && y_pointer == 46)
||(x_pointer == 95 && y_pointer == 46)
||(x_pointer == 96 && y_pointer == 46)
||(x_pointer == 97 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 99 && y_pointer == 46)
||(x_pointer == 100 && y_pointer == 46)
||(x_pointer == 101 && y_pointer == 46)
||(x_pointer == 102 && y_pointer == 46)
||(x_pointer == 103 && y_pointer == 46)
||(x_pointer == 104 && y_pointer == 46)
||(x_pointer == 105 && y_pointer == 46)
||(x_pointer == 106 && y_pointer == 46)
||(x_pointer == 107 && y_pointer == 46)
||(x_pointer == 108 && y_pointer == 46)
||(x_pointer == 109 && y_pointer == 46)
||(x_pointer == 110 && y_pointer == 46)
||(x_pointer == 111 && y_pointer == 46)
||(x_pointer == 112 && y_pointer == 46)
||(x_pointer == 113 && y_pointer == 46)
||(x_pointer == 114 && y_pointer == 46)
||(x_pointer == 115 && y_pointer == 46)
||(x_pointer == 116 && y_pointer == 46)
||(x_pointer == 117 && y_pointer == 46)
||(x_pointer == 118 && y_pointer == 46)
||(x_pointer == 119 && y_pointer == 46)
||(x_pointer == 120 && y_pointer == 46)
||(x_pointer == 121 && y_pointer == 46)
||(x_pointer == 122 && y_pointer == 46)
||(x_pointer == 123 && y_pointer == 46)
||(x_pointer == 124 && y_pointer == 46)
||(x_pointer == 125 && y_pointer == 46)
||(x_pointer == 126 && y_pointer == 46)
||(x_pointer == 127 && y_pointer == 46)
||(x_pointer == 128 && y_pointer == 46)
||(x_pointer == 129 && y_pointer == 46)
||(x_pointer == 130 && y_pointer == 46)
||(x_pointer == 131 && y_pointer == 46)
||(x_pointer == 132 && y_pointer == 46)
||(x_pointer == 133 && y_pointer == 46)
||(x_pointer == 134 && y_pointer == 46)
||(x_pointer == 135 && y_pointer == 46)
||(x_pointer == 136 && y_pointer == 46)
||(x_pointer == 137 && y_pointer == 46)
||(x_pointer == 138 && y_pointer == 46)
||(x_pointer == 139 && y_pointer == 46)
||(x_pointer == 140 && y_pointer == 46)
||(x_pointer == 141 && y_pointer == 46)
||(x_pointer == 142 && y_pointer == 46)
||(x_pointer == 143 && y_pointer == 46)
||(x_pointer == 144 && y_pointer == 46)
||(x_pointer == 145 && y_pointer == 46)
||(x_pointer == 146 && y_pointer == 46)
||(x_pointer == 147 && y_pointer == 46)
||(x_pointer == 148 && y_pointer == 46)
||(x_pointer == 149 && y_pointer == 46)
||(x_pointer == 150 && y_pointer == 46)
||(x_pointer == 151 && y_pointer == 46)
||(x_pointer == 152 && y_pointer == 46)
||(x_pointer == 153 && y_pointer == 46)
||(x_pointer == 154 && y_pointer == 46)
||(x_pointer == 32 && y_pointer == 47)
||(x_pointer == 33 && y_pointer == 47)
||(x_pointer == 34 && y_pointer == 47)
||(x_pointer == 35 && y_pointer == 47)
||(x_pointer == 36 && y_pointer == 47)
||(x_pointer == 37 && y_pointer == 47)
||(x_pointer == 38 && y_pointer == 47)
||(x_pointer == 39 && y_pointer == 47)
||(x_pointer == 40 && y_pointer == 47)
||(x_pointer == 32 && y_pointer == 48)
||(x_pointer == 33 && y_pointer == 48)
||(x_pointer == 34 && y_pointer == 48)
||(x_pointer == 35 && y_pointer == 48)
||(x_pointer == 36 && y_pointer == 48)
||(x_pointer == 37 && y_pointer == 48)
||(x_pointer == 38 && y_pointer == 48)
||(x_pointer == 39 && y_pointer == 48)
||(x_pointer == 40 && y_pointer == 48)
||(x_pointer == 32 && y_pointer == 49)
||(x_pointer == 33 && y_pointer == 49)
||(x_pointer == 34 && y_pointer == 49)
||(x_pointer == 35 && y_pointer == 49)
||(x_pointer == 36 && y_pointer == 49)
||(x_pointer == 37 && y_pointer == 49)
||(x_pointer == 38 && y_pointer == 49)
||(x_pointer == 39 && y_pointer == 49)
||(x_pointer == 40 && y_pointer == 49)
||(x_pointer == 32 && y_pointer == 50)
||(x_pointer == 33 && y_pointer == 50)
||(x_pointer == 34 && y_pointer == 50)
||(x_pointer == 35 && y_pointer == 50)
||(x_pointer == 36 && y_pointer == 50)
||(x_pointer == 37 && y_pointer == 50)
||(x_pointer == 38 && y_pointer == 50)
||(x_pointer == 39 && y_pointer == 50)
||(x_pointer == 40 && y_pointer == 50)
||(x_pointer == 32 && y_pointer == 51)
||(x_pointer == 33 && y_pointer == 51)
||(x_pointer == 34 && y_pointer == 51)
||(x_pointer == 35 && y_pointer == 51)
||(x_pointer == 36 && y_pointer == 51)
||(x_pointer == 37 && y_pointer == 51)
||(x_pointer == 38 && y_pointer == 51)
||(x_pointer == 39 && y_pointer == 51)
||(x_pointer == 40 && y_pointer == 51)
||(x_pointer == 32 && y_pointer == 52)
||(x_pointer == 33 && y_pointer == 52)
||(x_pointer == 34 && y_pointer == 52)
||(x_pointer == 35 && y_pointer == 52)
||(x_pointer == 36 && y_pointer == 52)
||(x_pointer == 37 && y_pointer == 52)
||(x_pointer == 38 && y_pointer == 52)
||(x_pointer == 39 && y_pointer == 52)
||(x_pointer == 40 && y_pointer == 52)
||(x_pointer == 32 && y_pointer == 53)
||(x_pointer == 33 && y_pointer == 53)
||(x_pointer == 34 && y_pointer == 53)
||(x_pointer == 35 && y_pointer == 53)
||(x_pointer == 36 && y_pointer == 53)
||(x_pointer == 37 && y_pointer == 53)
||(x_pointer == 38 && y_pointer == 53)
||(x_pointer == 39 && y_pointer == 53)
||(x_pointer == 40 && y_pointer == 53)
||(x_pointer == 32 && y_pointer == 54)
||(x_pointer == 33 && y_pointer == 54)
||(x_pointer == 34 && y_pointer == 54)
||(x_pointer == 35 && y_pointer == 54)
||(x_pointer == 36 && y_pointer == 54)
||(x_pointer == 37 && y_pointer == 54)
||(x_pointer == 38 && y_pointer == 54)
||(x_pointer == 39 && y_pointer == 54)
||(x_pointer == 40 && y_pointer == 54)
||(x_pointer == 32 && y_pointer == 55)
||(x_pointer == 33 && y_pointer == 55)
||(x_pointer == 34 && y_pointer == 55)
||(x_pointer == 35 && y_pointer == 55)
||(x_pointer == 36 && y_pointer == 55)
||(x_pointer == 37 && y_pointer == 55)
||(x_pointer == 38 && y_pointer == 55)
||(x_pointer == 39 && y_pointer == 55)
||(x_pointer == 40 && y_pointer == 55)
||(x_pointer == 32 && y_pointer == 56)
||(x_pointer == 33 && y_pointer == 56)
||(x_pointer == 34 && y_pointer == 56)
||(x_pointer == 35 && y_pointer == 56)
||(x_pointer == 36 && y_pointer == 56)
||(x_pointer == 37 && y_pointer == 56)
||(x_pointer == 38 && y_pointer == 56)
||(x_pointer == 39 && y_pointer == 56)
||(x_pointer == 40 && y_pointer == 56)
||(x_pointer == 32 && y_pointer == 57)
||(x_pointer == 33 && y_pointer == 57)
||(x_pointer == 34 && y_pointer == 57)
||(x_pointer == 35 && y_pointer == 57)
||(x_pointer == 36 && y_pointer == 57)
||(x_pointer == 37 && y_pointer == 57)
||(x_pointer == 38 && y_pointer == 57)
||(x_pointer == 39 && y_pointer == 57)
||(x_pointer == 40 && y_pointer == 57)
||(x_pointer == 32 && y_pointer == 58)
||(x_pointer == 33 && y_pointer == 58)
||(x_pointer == 34 && y_pointer == 58)
||(x_pointer == 35 && y_pointer == 58)
||(x_pointer == 36 && y_pointer == 58)
||(x_pointer == 37 && y_pointer == 58)
||(x_pointer == 38 && y_pointer == 58)
||(x_pointer == 39 && y_pointer == 58)
||(x_pointer == 40 && y_pointer == 58)
||(x_pointer == 32 && y_pointer == 59)
||(x_pointer == 33 && y_pointer == 59)
||(x_pointer == 34 && y_pointer == 59)
||(x_pointer == 35 && y_pointer == 59)
||(x_pointer == 36 && y_pointer == 59)
||(x_pointer == 37 && y_pointer == 59)
||(x_pointer == 38 && y_pointer == 59)
||(x_pointer == 39 && y_pointer == 59)
||(x_pointer == 40 && y_pointer == 59)
||(x_pointer == 32 && y_pointer == 60)
||(x_pointer == 33 && y_pointer == 60)
||(x_pointer == 34 && y_pointer == 60)
||(x_pointer == 35 && y_pointer == 60)
||(x_pointer == 36 && y_pointer == 60)
||(x_pointer == 37 && y_pointer == 60)
||(x_pointer == 38 && y_pointer == 60)
||(x_pointer == 39 && y_pointer == 60)
||(x_pointer == 40 && y_pointer == 60)
||(x_pointer == 32 && y_pointer == 61)
||(x_pointer == 33 && y_pointer == 61)
||(x_pointer == 34 && y_pointer == 61)
||(x_pointer == 35 && y_pointer == 61)
||(x_pointer == 36 && y_pointer == 61)
||(x_pointer == 37 && y_pointer == 61)
||(x_pointer == 38 && y_pointer == 61)
||(x_pointer == 39 && y_pointer == 61)
||(x_pointer == 40 && y_pointer == 61)
||(x_pointer == 32 && y_pointer == 62)
||(x_pointer == 33 && y_pointer == 62)
||(x_pointer == 34 && y_pointer == 62)
||(x_pointer == 35 && y_pointer == 62)
||(x_pointer == 36 && y_pointer == 62)
||(x_pointer == 37 && y_pointer == 62)
||(x_pointer == 38 && y_pointer == 62)
||(x_pointer == 39 && y_pointer == 62)
||(x_pointer == 40 && y_pointer == 62)
||(x_pointer == 68 && y_pointer == 62)
||(x_pointer == 69 && y_pointer == 62)
||(x_pointer == 70 && y_pointer == 62)
||(x_pointer == 71 && y_pointer == 62)
||(x_pointer == 72 && y_pointer == 62)
||(x_pointer == 73 && y_pointer == 62)
||(x_pointer == 74 && y_pointer == 62)
||(x_pointer == 75 && y_pointer == 62)
||(x_pointer == 76 && y_pointer == 62)
||(x_pointer == 77 && y_pointer == 62)
||(x_pointer == 78 && y_pointer == 62)
||(x_pointer == 79 && y_pointer == 62)
||(x_pointer == 80 && y_pointer == 62)
||(x_pointer == 81 && y_pointer == 62)
||(x_pointer == 82 && y_pointer == 62)
||(x_pointer == 83 && y_pointer == 62)
||(x_pointer == 84 && y_pointer == 62)
||(x_pointer == 32 && y_pointer == 63)
||(x_pointer == 33 && y_pointer == 63)
||(x_pointer == 34 && y_pointer == 63)
||(x_pointer == 35 && y_pointer == 63)
||(x_pointer == 36 && y_pointer == 63)
||(x_pointer == 37 && y_pointer == 63)
||(x_pointer == 38 && y_pointer == 63)
||(x_pointer == 39 && y_pointer == 63)
||(x_pointer == 40 && y_pointer == 63)
||(x_pointer == 68 && y_pointer == 63)
||(x_pointer == 69 && y_pointer == 63)
||(x_pointer == 70 && y_pointer == 63)
||(x_pointer == 71 && y_pointer == 63)
||(x_pointer == 72 && y_pointer == 63)
||(x_pointer == 73 && y_pointer == 63)
||(x_pointer == 74 && y_pointer == 63)
||(x_pointer == 75 && y_pointer == 63)
||(x_pointer == 76 && y_pointer == 63)
||(x_pointer == 77 && y_pointer == 63)
||(x_pointer == 78 && y_pointer == 63)
||(x_pointer == 79 && y_pointer == 63)
||(x_pointer == 80 && y_pointer == 63)
||(x_pointer == 81 && y_pointer == 63)
||(x_pointer == 82 && y_pointer == 63)
||(x_pointer == 83 && y_pointer == 63)
||(x_pointer == 84 && y_pointer == 63)
||(x_pointer == 32 && y_pointer == 64)
||(x_pointer == 33 && y_pointer == 64)
||(x_pointer == 34 && y_pointer == 64)
||(x_pointer == 35 && y_pointer == 64)
||(x_pointer == 36 && y_pointer == 64)
||(x_pointer == 37 && y_pointer == 64)
||(x_pointer == 38 && y_pointer == 64)
||(x_pointer == 39 && y_pointer == 64)
||(x_pointer == 40 && y_pointer == 64)
||(x_pointer == 68 && y_pointer == 64)
||(x_pointer == 69 && y_pointer == 64)
||(x_pointer == 70 && y_pointer == 64)
||(x_pointer == 71 && y_pointer == 64)
||(x_pointer == 72 && y_pointer == 64)
||(x_pointer == 73 && y_pointer == 64)
||(x_pointer == 74 && y_pointer == 64)
||(x_pointer == 75 && y_pointer == 64)
||(x_pointer == 76 && y_pointer == 64)
||(x_pointer == 77 && y_pointer == 64)
||(x_pointer == 78 && y_pointer == 64)
||(x_pointer == 79 && y_pointer == 64)
||(x_pointer == 80 && y_pointer == 64)
||(x_pointer == 81 && y_pointer == 64)
||(x_pointer == 82 && y_pointer == 64)
||(x_pointer == 83 && y_pointer == 64)
||(x_pointer == 84 && y_pointer == 64)
||(x_pointer == 32 && y_pointer == 65)
||(x_pointer == 33 && y_pointer == 65)
||(x_pointer == 34 && y_pointer == 65)
||(x_pointer == 35 && y_pointer == 65)
||(x_pointer == 36 && y_pointer == 65)
||(x_pointer == 37 && y_pointer == 65)
||(x_pointer == 38 && y_pointer == 65)
||(x_pointer == 39 && y_pointer == 65)
||(x_pointer == 40 && y_pointer == 65)
||(x_pointer == 68 && y_pointer == 65)
||(x_pointer == 69 && y_pointer == 65)
||(x_pointer == 70 && y_pointer == 65)
||(x_pointer == 71 && y_pointer == 65)
||(x_pointer == 72 && y_pointer == 65)
||(x_pointer == 73 && y_pointer == 65)
||(x_pointer == 74 && y_pointer == 65)
||(x_pointer == 75 && y_pointer == 65)
||(x_pointer == 76 && y_pointer == 65)
||(x_pointer == 77 && y_pointer == 65)
||(x_pointer == 78 && y_pointer == 65)
||(x_pointer == 79 && y_pointer == 65)
||(x_pointer == 80 && y_pointer == 65)
||(x_pointer == 81 && y_pointer == 65)
||(x_pointer == 82 && y_pointer == 65)
||(x_pointer == 83 && y_pointer == 65)
||(x_pointer == 84 && y_pointer == 65)
||(x_pointer == 32 && y_pointer == 66)
||(x_pointer == 33 && y_pointer == 66)
||(x_pointer == 34 && y_pointer == 66)
||(x_pointer == 35 && y_pointer == 66)
||(x_pointer == 36 && y_pointer == 66)
||(x_pointer == 37 && y_pointer == 66)
||(x_pointer == 38 && y_pointer == 66)
||(x_pointer == 39 && y_pointer == 66)
||(x_pointer == 40 && y_pointer == 66)
||(x_pointer == 68 && y_pointer == 66)
||(x_pointer == 69 && y_pointer == 66)
||(x_pointer == 70 && y_pointer == 66)
||(x_pointer == 71 && y_pointer == 66)
||(x_pointer == 72 && y_pointer == 66)
||(x_pointer == 73 && y_pointer == 66)
||(x_pointer == 74 && y_pointer == 66)
||(x_pointer == 75 && y_pointer == 66)
||(x_pointer == 76 && y_pointer == 66)
||(x_pointer == 77 && y_pointer == 66)
||(x_pointer == 78 && y_pointer == 66)
||(x_pointer == 79 && y_pointer == 66)
||(x_pointer == 80 && y_pointer == 66)
||(x_pointer == 81 && y_pointer == 66)
||(x_pointer == 82 && y_pointer == 66)
||(x_pointer == 83 && y_pointer == 66)
||(x_pointer == 84 && y_pointer == 66)
||(x_pointer == 32 && y_pointer == 67)
||(x_pointer == 33 && y_pointer == 67)
||(x_pointer == 34 && y_pointer == 67)
||(x_pointer == 35 && y_pointer == 67)
||(x_pointer == 36 && y_pointer == 67)
||(x_pointer == 37 && y_pointer == 67)
||(x_pointer == 38 && y_pointer == 67)
||(x_pointer == 39 && y_pointer == 67)
||(x_pointer == 40 && y_pointer == 67)
||(x_pointer == 68 && y_pointer == 67)
||(x_pointer == 69 && y_pointer == 67)
||(x_pointer == 70 && y_pointer == 67)
||(x_pointer == 71 && y_pointer == 67)
||(x_pointer == 72 && y_pointer == 67)
||(x_pointer == 73 && y_pointer == 67)
||(x_pointer == 74 && y_pointer == 67)
||(x_pointer == 75 && y_pointer == 67)
||(x_pointer == 76 && y_pointer == 67)
||(x_pointer == 77 && y_pointer == 67)
||(x_pointer == 78 && y_pointer == 67)
||(x_pointer == 79 && y_pointer == 67)
||(x_pointer == 80 && y_pointer == 67)
||(x_pointer == 81 && y_pointer == 67)
||(x_pointer == 82 && y_pointer == 67)
||(x_pointer == 83 && y_pointer == 67)
||(x_pointer == 84 && y_pointer == 67)
||(x_pointer == 68 && y_pointer == 68)
||(x_pointer == 69 && y_pointer == 68)
||(x_pointer == 70 && y_pointer == 68)
||(x_pointer == 71 && y_pointer == 68)
||(x_pointer == 72 && y_pointer == 68)
||(x_pointer == 73 && y_pointer == 68)
||(x_pointer == 74 && y_pointer == 68)
||(x_pointer == 75 && y_pointer == 68)
||(x_pointer == 76 && y_pointer == 68)
||(x_pointer == 77 && y_pointer == 68)
||(x_pointer == 78 && y_pointer == 68)
||(x_pointer == 79 && y_pointer == 68)
||(x_pointer == 80 && y_pointer == 68)
||(x_pointer == 81 && y_pointer == 68)
||(x_pointer == 82 && y_pointer == 68)
||(x_pointer == 83 && y_pointer == 68)
||(x_pointer == 84 && y_pointer == 68)
||(x_pointer == 110 && y_pointer == 68)
||(x_pointer == 111 && y_pointer == 68)
||(x_pointer == 112 && y_pointer == 68)
||(x_pointer == 113 && y_pointer == 68)
||(x_pointer == 114 && y_pointer == 68)
||(x_pointer == 115 && y_pointer == 68)
||(x_pointer == 116 && y_pointer == 68)
||(x_pointer == 117 && y_pointer == 68)
||(x_pointer == 118 && y_pointer == 68)
||(x_pointer == 68 && y_pointer == 69)
||(x_pointer == 69 && y_pointer == 69)
||(x_pointer == 70 && y_pointer == 69)
||(x_pointer == 71 && y_pointer == 69)
||(x_pointer == 72 && y_pointer == 69)
||(x_pointer == 73 && y_pointer == 69)
||(x_pointer == 74 && y_pointer == 69)
||(x_pointer == 75 && y_pointer == 69)
||(x_pointer == 76 && y_pointer == 69)
||(x_pointer == 77 && y_pointer == 69)
||(x_pointer == 78 && y_pointer == 69)
||(x_pointer == 79 && y_pointer == 69)
||(x_pointer == 80 && y_pointer == 69)
||(x_pointer == 81 && y_pointer == 69)
||(x_pointer == 82 && y_pointer == 69)
||(x_pointer == 83 && y_pointer == 69)
||(x_pointer == 84 && y_pointer == 69)
||(x_pointer == 110 && y_pointer == 69)
||(x_pointer == 111 && y_pointer == 69)
||(x_pointer == 112 && y_pointer == 69)
||(x_pointer == 113 && y_pointer == 69)
||(x_pointer == 114 && y_pointer == 69)
||(x_pointer == 115 && y_pointer == 69)
||(x_pointer == 116 && y_pointer == 69)
||(x_pointer == 117 && y_pointer == 69)
||(x_pointer == 118 && y_pointer == 69)
||(x_pointer == 68 && y_pointer == 70)
||(x_pointer == 69 && y_pointer == 70)
||(x_pointer == 70 && y_pointer == 70)
||(x_pointer == 71 && y_pointer == 70)
||(x_pointer == 72 && y_pointer == 70)
||(x_pointer == 73 && y_pointer == 70)
||(x_pointer == 74 && y_pointer == 70)
||(x_pointer == 75 && y_pointer == 70)
||(x_pointer == 76 && y_pointer == 70)
||(x_pointer == 77 && y_pointer == 70)
||(x_pointer == 78 && y_pointer == 70)
||(x_pointer == 79 && y_pointer == 70)
||(x_pointer == 80 && y_pointer == 70)
||(x_pointer == 81 && y_pointer == 70)
||(x_pointer == 82 && y_pointer == 70)
||(x_pointer == 83 && y_pointer == 70)
||(x_pointer == 84 && y_pointer == 70)
||(x_pointer == 110 && y_pointer == 70)
||(x_pointer == 111 && y_pointer == 70)
||(x_pointer == 112 && y_pointer == 70)
||(x_pointer == 113 && y_pointer == 70)
||(x_pointer == 114 && y_pointer == 70)
||(x_pointer == 115 && y_pointer == 70)
||(x_pointer == 116 && y_pointer == 70)
||(x_pointer == 117 && y_pointer == 70)
||(x_pointer == 118 && y_pointer == 70)
||(x_pointer == 68 && y_pointer == 71)
||(x_pointer == 69 && y_pointer == 71)
||(x_pointer == 70 && y_pointer == 71)
||(x_pointer == 71 && y_pointer == 71)
||(x_pointer == 72 && y_pointer == 71)
||(x_pointer == 73 && y_pointer == 71)
||(x_pointer == 74 && y_pointer == 71)
||(x_pointer == 75 && y_pointer == 71)
||(x_pointer == 76 && y_pointer == 71)
||(x_pointer == 77 && y_pointer == 71)
||(x_pointer == 78 && y_pointer == 71)
||(x_pointer == 79 && y_pointer == 71)
||(x_pointer == 80 && y_pointer == 71)
||(x_pointer == 81 && y_pointer == 71)
||(x_pointer == 82 && y_pointer == 71)
||(x_pointer == 83 && y_pointer == 71)
||(x_pointer == 84 && y_pointer == 71)
||(x_pointer == 110 && y_pointer == 71)
||(x_pointer == 111 && y_pointer == 71)
||(x_pointer == 112 && y_pointer == 71)
||(x_pointer == 113 && y_pointer == 71)
||(x_pointer == 114 && y_pointer == 71)
||(x_pointer == 115 && y_pointer == 71)
||(x_pointer == 116 && y_pointer == 71)
||(x_pointer == 117 && y_pointer == 71)
||(x_pointer == 118 && y_pointer == 71)
||(x_pointer == 68 && y_pointer == 72)
||(x_pointer == 69 && y_pointer == 72)
||(x_pointer == 70 && y_pointer == 72)
||(x_pointer == 71 && y_pointer == 72)
||(x_pointer == 72 && y_pointer == 72)
||(x_pointer == 73 && y_pointer == 72)
||(x_pointer == 74 && y_pointer == 72)
||(x_pointer == 75 && y_pointer == 72)
||(x_pointer == 76 && y_pointer == 72)
||(x_pointer == 77 && y_pointer == 72)
||(x_pointer == 78 && y_pointer == 72)
||(x_pointer == 79 && y_pointer == 72)
||(x_pointer == 80 && y_pointer == 72)
||(x_pointer == 81 && y_pointer == 72)
||(x_pointer == 82 && y_pointer == 72)
||(x_pointer == 83 && y_pointer == 72)
||(x_pointer == 84 && y_pointer == 72)
||(x_pointer == 110 && y_pointer == 72)
||(x_pointer == 111 && y_pointer == 72)
||(x_pointer == 112 && y_pointer == 72)
||(x_pointer == 113 && y_pointer == 72)
||(x_pointer == 114 && y_pointer == 72)
||(x_pointer == 115 && y_pointer == 72)
||(x_pointer == 116 && y_pointer == 72)
||(x_pointer == 117 && y_pointer == 72)
||(x_pointer == 118 && y_pointer == 72)
||(x_pointer == 68 && y_pointer == 73)
||(x_pointer == 69 && y_pointer == 73)
||(x_pointer == 70 && y_pointer == 73)
||(x_pointer == 71 && y_pointer == 73)
||(x_pointer == 72 && y_pointer == 73)
||(x_pointer == 73 && y_pointer == 73)
||(x_pointer == 74 && y_pointer == 73)
||(x_pointer == 75 && y_pointer == 73)
||(x_pointer == 76 && y_pointer == 73)
||(x_pointer == 77 && y_pointer == 73)
||(x_pointer == 78 && y_pointer == 73)
||(x_pointer == 79 && y_pointer == 73)
||(x_pointer == 80 && y_pointer == 73)
||(x_pointer == 81 && y_pointer == 73)
||(x_pointer == 82 && y_pointer == 73)
||(x_pointer == 83 && y_pointer == 73)
||(x_pointer == 84 && y_pointer == 73)
||(x_pointer == 110 && y_pointer == 73)
||(x_pointer == 111 && y_pointer == 73)
||(x_pointer == 112 && y_pointer == 73)
||(x_pointer == 113 && y_pointer == 73)
||(x_pointer == 114 && y_pointer == 73)
||(x_pointer == 115 && y_pointer == 73)
||(x_pointer == 116 && y_pointer == 73)
||(x_pointer == 117 && y_pointer == 73)
||(x_pointer == 118 && y_pointer == 73)
||(x_pointer == 68 && y_pointer == 74)
||(x_pointer == 69 && y_pointer == 74)
||(x_pointer == 70 && y_pointer == 74)
||(x_pointer == 71 && y_pointer == 74)
||(x_pointer == 72 && y_pointer == 74)
||(x_pointer == 73 && y_pointer == 74)
||(x_pointer == 74 && y_pointer == 74)
||(x_pointer == 75 && y_pointer == 74)
||(x_pointer == 76 && y_pointer == 74)
||(x_pointer == 77 && y_pointer == 74)
||(x_pointer == 78 && y_pointer == 74)
||(x_pointer == 79 && y_pointer == 74)
||(x_pointer == 80 && y_pointer == 74)
||(x_pointer == 81 && y_pointer == 74)
||(x_pointer == 82 && y_pointer == 74)
||(x_pointer == 83 && y_pointer == 74)
||(x_pointer == 84 && y_pointer == 74)
||(x_pointer == 110 && y_pointer == 74)
||(x_pointer == 111 && y_pointer == 74)
||(x_pointer == 112 && y_pointer == 74)
||(x_pointer == 113 && y_pointer == 74)
||(x_pointer == 114 && y_pointer == 74)
||(x_pointer == 115 && y_pointer == 74)
||(x_pointer == 116 && y_pointer == 74)
||(x_pointer == 117 && y_pointer == 74)
||(x_pointer == 118 && y_pointer == 74)
||(x_pointer == 68 && y_pointer == 75)
||(x_pointer == 69 && y_pointer == 75)
||(x_pointer == 70 && y_pointer == 75)
||(x_pointer == 71 && y_pointer == 75)
||(x_pointer == 72 && y_pointer == 75)
||(x_pointer == 73 && y_pointer == 75)
||(x_pointer == 74 && y_pointer == 75)
||(x_pointer == 75 && y_pointer == 75)
||(x_pointer == 76 && y_pointer == 75)
||(x_pointer == 77 && y_pointer == 75)
||(x_pointer == 78 && y_pointer == 75)
||(x_pointer == 79 && y_pointer == 75)
||(x_pointer == 80 && y_pointer == 75)
||(x_pointer == 81 && y_pointer == 75)
||(x_pointer == 82 && y_pointer == 75)
||(x_pointer == 83 && y_pointer == 75)
||(x_pointer == 84 && y_pointer == 75)
||(x_pointer == 110 && y_pointer == 75)
||(x_pointer == 111 && y_pointer == 75)
||(x_pointer == 112 && y_pointer == 75)
||(x_pointer == 113 && y_pointer == 75)
||(x_pointer == 114 && y_pointer == 75)
||(x_pointer == 115 && y_pointer == 75)
||(x_pointer == 116 && y_pointer == 75)
||(x_pointer == 117 && y_pointer == 75)
||(x_pointer == 118 && y_pointer == 75)
||(x_pointer == 68 && y_pointer == 76)
||(x_pointer == 69 && y_pointer == 76)
||(x_pointer == 70 && y_pointer == 76)
||(x_pointer == 71 && y_pointer == 76)
||(x_pointer == 72 && y_pointer == 76)
||(x_pointer == 73 && y_pointer == 76)
||(x_pointer == 74 && y_pointer == 76)
||(x_pointer == 75 && y_pointer == 76)
||(x_pointer == 76 && y_pointer == 76)
||(x_pointer == 77 && y_pointer == 76)
||(x_pointer == 78 && y_pointer == 76)
||(x_pointer == 79 && y_pointer == 76)
||(x_pointer == 80 && y_pointer == 76)
||(x_pointer == 81 && y_pointer == 76)
||(x_pointer == 82 && y_pointer == 76)
||(x_pointer == 83 && y_pointer == 76)
||(x_pointer == 84 && y_pointer == 76)
||(x_pointer == 110 && y_pointer == 76)
||(x_pointer == 111 && y_pointer == 76)
||(x_pointer == 112 && y_pointer == 76)
||(x_pointer == 113 && y_pointer == 76)
||(x_pointer == 114 && y_pointer == 76)
||(x_pointer == 115 && y_pointer == 76)
||(x_pointer == 116 && y_pointer == 76)
||(x_pointer == 117 && y_pointer == 76)
||(x_pointer == 118 && y_pointer == 76)
||(x_pointer == 110 && y_pointer == 77)
||(x_pointer == 111 && y_pointer == 77)
||(x_pointer == 112 && y_pointer == 77)
||(x_pointer == 113 && y_pointer == 77)
||(x_pointer == 114 && y_pointer == 77)
||(x_pointer == 115 && y_pointer == 77)
||(x_pointer == 116 && y_pointer == 77)
||(x_pointer == 117 && y_pointer == 77)
||(x_pointer == 118 && y_pointer == 77)
||(x_pointer == 110 && y_pointer == 78)
||(x_pointer == 111 && y_pointer == 78)
||(x_pointer == 112 && y_pointer == 78)
||(x_pointer == 113 && y_pointer == 78)
||(x_pointer == 114 && y_pointer == 78)
||(x_pointer == 115 && y_pointer == 78)
||(x_pointer == 116 && y_pointer == 78)
||(x_pointer == 117 && y_pointer == 78)
||(x_pointer == 118 && y_pointer == 78)
||(x_pointer == 110 && y_pointer == 79)
||(x_pointer == 111 && y_pointer == 79)
||(x_pointer == 112 && y_pointer == 79)
||(x_pointer == 113 && y_pointer == 79)
||(x_pointer == 114 && y_pointer == 79)
||(x_pointer == 115 && y_pointer == 79)
||(x_pointer == 116 && y_pointer == 79)
||(x_pointer == 117 && y_pointer == 79)
||(x_pointer == 118 && y_pointer == 79)
||(x_pointer == 110 && y_pointer == 80)
||(x_pointer == 111 && y_pointer == 80)
||(x_pointer == 112 && y_pointer == 80)
||(x_pointer == 113 && y_pointer == 80)
||(x_pointer == 114 && y_pointer == 80)
||(x_pointer == 115 && y_pointer == 80)
||(x_pointer == 116 && y_pointer == 80)
||(x_pointer == 117 && y_pointer == 80)
||(x_pointer == 118 && y_pointer == 80)
||(x_pointer == 110 && y_pointer == 81)
||(x_pointer == 111 && y_pointer == 81)
||(x_pointer == 112 && y_pointer == 81)
||(x_pointer == 113 && y_pointer == 81)
||(x_pointer == 114 && y_pointer == 81)
||(x_pointer == 115 && y_pointer == 81)
||(x_pointer == 116 && y_pointer == 81)
||(x_pointer == 117 && y_pointer == 81)
||(x_pointer == 118 && y_pointer == 81)
||(x_pointer == 110 && y_pointer == 82)
||(x_pointer == 111 && y_pointer == 82)
||(x_pointer == 112 && y_pointer == 82)
||(x_pointer == 113 && y_pointer == 82)
||(x_pointer == 114 && y_pointer == 82)
||(x_pointer == 115 && y_pointer == 82)
||(x_pointer == 116 && y_pointer == 82)
||(x_pointer == 117 && y_pointer == 82)
||(x_pointer == 118 && y_pointer == 82)
||(x_pointer == 5 && y_pointer == 83)
||(x_pointer == 6 && y_pointer == 83)
||(x_pointer == 7 && y_pointer == 83)
||(x_pointer == 8 && y_pointer == 83)
||(x_pointer == 9 && y_pointer == 83)
||(x_pointer == 10 && y_pointer == 83)
||(x_pointer == 11 && y_pointer == 83)
||(x_pointer == 12 && y_pointer == 83)
||(x_pointer == 13 && y_pointer == 83)
||(x_pointer == 14 && y_pointer == 83)
||(x_pointer == 15 && y_pointer == 83)
||(x_pointer == 16 && y_pointer == 83)
||(x_pointer == 17 && y_pointer == 83)
||(x_pointer == 18 && y_pointer == 83)
||(x_pointer == 19 && y_pointer == 83)
||(x_pointer == 20 && y_pointer == 83)
||(x_pointer == 21 && y_pointer == 83)
||(x_pointer == 22 && y_pointer == 83)
||(x_pointer == 23 && y_pointer == 83)
||(x_pointer == 24 && y_pointer == 83)
||(x_pointer == 25 && y_pointer == 83)
||(x_pointer == 26 && y_pointer == 83)
||(x_pointer == 27 && y_pointer == 83)
||(x_pointer == 28 && y_pointer == 83)
||(x_pointer == 29 && y_pointer == 83)
||(x_pointer == 30 && y_pointer == 83)
||(x_pointer == 31 && y_pointer == 83)
||(x_pointer == 32 && y_pointer == 83)
||(x_pointer == 33 && y_pointer == 83)
||(x_pointer == 34 && y_pointer == 83)
||(x_pointer == 35 && y_pointer == 83)
||(x_pointer == 36 && y_pointer == 83)
||(x_pointer == 37 && y_pointer == 83)
||(x_pointer == 38 && y_pointer == 83)
||(x_pointer == 39 && y_pointer == 83)
||(x_pointer == 40 && y_pointer == 83)
||(x_pointer == 41 && y_pointer == 83)
||(x_pointer == 42 && y_pointer == 83)
||(x_pointer == 43 && y_pointer == 83)
||(x_pointer == 44 && y_pointer == 83)
||(x_pointer == 45 && y_pointer == 83)
||(x_pointer == 46 && y_pointer == 83)
||(x_pointer == 47 && y_pointer == 83)
||(x_pointer == 48 && y_pointer == 83)
||(x_pointer == 49 && y_pointer == 83)
||(x_pointer == 50 && y_pointer == 83)
||(x_pointer == 51 && y_pointer == 83)
||(x_pointer == 52 && y_pointer == 83)
||(x_pointer == 53 && y_pointer == 83)
||(x_pointer == 54 && y_pointer == 83)
||(x_pointer == 55 && y_pointer == 83)
||(x_pointer == 56 && y_pointer == 83)
||(x_pointer == 57 && y_pointer == 83)
||(x_pointer == 58 && y_pointer == 83)
||(x_pointer == 110 && y_pointer == 83)
||(x_pointer == 111 && y_pointer == 83)
||(x_pointer == 112 && y_pointer == 83)
||(x_pointer == 113 && y_pointer == 83)
||(x_pointer == 114 && y_pointer == 83)
||(x_pointer == 115 && y_pointer == 83)
||(x_pointer == 116 && y_pointer == 83)
||(x_pointer == 117 && y_pointer == 83)
||(x_pointer == 118 && y_pointer == 83)
||(x_pointer == 5 && y_pointer == 84)
||(x_pointer == 6 && y_pointer == 84)
||(x_pointer == 7 && y_pointer == 84)
||(x_pointer == 8 && y_pointer == 84)
||(x_pointer == 9 && y_pointer == 84)
||(x_pointer == 10 && y_pointer == 84)
||(x_pointer == 11 && y_pointer == 84)
||(x_pointer == 12 && y_pointer == 84)
||(x_pointer == 13 && y_pointer == 84)
||(x_pointer == 14 && y_pointer == 84)
||(x_pointer == 15 && y_pointer == 84)
||(x_pointer == 16 && y_pointer == 84)
||(x_pointer == 17 && y_pointer == 84)
||(x_pointer == 18 && y_pointer == 84)
||(x_pointer == 19 && y_pointer == 84)
||(x_pointer == 20 && y_pointer == 84)
||(x_pointer == 21 && y_pointer == 84)
||(x_pointer == 22 && y_pointer == 84)
||(x_pointer == 23 && y_pointer == 84)
||(x_pointer == 24 && y_pointer == 84)
||(x_pointer == 25 && y_pointer == 84)
||(x_pointer == 26 && y_pointer == 84)
||(x_pointer == 27 && y_pointer == 84)
||(x_pointer == 28 && y_pointer == 84)
||(x_pointer == 29 && y_pointer == 84)
||(x_pointer == 30 && y_pointer == 84)
||(x_pointer == 31 && y_pointer == 84)
||(x_pointer == 32 && y_pointer == 84)
||(x_pointer == 33 && y_pointer == 84)
||(x_pointer == 34 && y_pointer == 84)
||(x_pointer == 35 && y_pointer == 84)
||(x_pointer == 36 && y_pointer == 84)
||(x_pointer == 37 && y_pointer == 84)
||(x_pointer == 38 && y_pointer == 84)
||(x_pointer == 39 && y_pointer == 84)
||(x_pointer == 40 && y_pointer == 84)
||(x_pointer == 41 && y_pointer == 84)
||(x_pointer == 42 && y_pointer == 84)
||(x_pointer == 43 && y_pointer == 84)
||(x_pointer == 44 && y_pointer == 84)
||(x_pointer == 45 && y_pointer == 84)
||(x_pointer == 46 && y_pointer == 84)
||(x_pointer == 47 && y_pointer == 84)
||(x_pointer == 48 && y_pointer == 84)
||(x_pointer == 49 && y_pointer == 84)
||(x_pointer == 50 && y_pointer == 84)
||(x_pointer == 51 && y_pointer == 84)
||(x_pointer == 52 && y_pointer == 84)
||(x_pointer == 53 && y_pointer == 84)
||(x_pointer == 54 && y_pointer == 84)
||(x_pointer == 55 && y_pointer == 84)
||(x_pointer == 56 && y_pointer == 84)
||(x_pointer == 57 && y_pointer == 84)
||(x_pointer == 58 && y_pointer == 84)
||(x_pointer == 110 && y_pointer == 84)
||(x_pointer == 111 && y_pointer == 84)
||(x_pointer == 112 && y_pointer == 84)
||(x_pointer == 113 && y_pointer == 84)
||(x_pointer == 114 && y_pointer == 84)
||(x_pointer == 115 && y_pointer == 84)
||(x_pointer == 116 && y_pointer == 84)
||(x_pointer == 117 && y_pointer == 84)
||(x_pointer == 118 && y_pointer == 84)
||(x_pointer == 5 && y_pointer == 85)
||(x_pointer == 6 && y_pointer == 85)
||(x_pointer == 7 && y_pointer == 85)
||(x_pointer == 8 && y_pointer == 85)
||(x_pointer == 9 && y_pointer == 85)
||(x_pointer == 10 && y_pointer == 85)
||(x_pointer == 11 && y_pointer == 85)
||(x_pointer == 12 && y_pointer == 85)
||(x_pointer == 13 && y_pointer == 85)
||(x_pointer == 14 && y_pointer == 85)
||(x_pointer == 15 && y_pointer == 85)
||(x_pointer == 16 && y_pointer == 85)
||(x_pointer == 17 && y_pointer == 85)
||(x_pointer == 18 && y_pointer == 85)
||(x_pointer == 19 && y_pointer == 85)
||(x_pointer == 20 && y_pointer == 85)
||(x_pointer == 21 && y_pointer == 85)
||(x_pointer == 22 && y_pointer == 85)
||(x_pointer == 23 && y_pointer == 85)
||(x_pointer == 24 && y_pointer == 85)
||(x_pointer == 25 && y_pointer == 85)
||(x_pointer == 26 && y_pointer == 85)
||(x_pointer == 27 && y_pointer == 85)
||(x_pointer == 28 && y_pointer == 85)
||(x_pointer == 29 && y_pointer == 85)
||(x_pointer == 30 && y_pointer == 85)
||(x_pointer == 31 && y_pointer == 85)
||(x_pointer == 32 && y_pointer == 85)
||(x_pointer == 33 && y_pointer == 85)
||(x_pointer == 34 && y_pointer == 85)
||(x_pointer == 35 && y_pointer == 85)
||(x_pointer == 36 && y_pointer == 85)
||(x_pointer == 37 && y_pointer == 85)
||(x_pointer == 38 && y_pointer == 85)
||(x_pointer == 39 && y_pointer == 85)
||(x_pointer == 40 && y_pointer == 85)
||(x_pointer == 41 && y_pointer == 85)
||(x_pointer == 42 && y_pointer == 85)
||(x_pointer == 43 && y_pointer == 85)
||(x_pointer == 44 && y_pointer == 85)
||(x_pointer == 45 && y_pointer == 85)
||(x_pointer == 46 && y_pointer == 85)
||(x_pointer == 47 && y_pointer == 85)
||(x_pointer == 48 && y_pointer == 85)
||(x_pointer == 49 && y_pointer == 85)
||(x_pointer == 50 && y_pointer == 85)
||(x_pointer == 51 && y_pointer == 85)
||(x_pointer == 52 && y_pointer == 85)
||(x_pointer == 53 && y_pointer == 85)
||(x_pointer == 54 && y_pointer == 85)
||(x_pointer == 55 && y_pointer == 85)
||(x_pointer == 56 && y_pointer == 85)
||(x_pointer == 57 && y_pointer == 85)
||(x_pointer == 58 && y_pointer == 85)
||(x_pointer == 110 && y_pointer == 85)
||(x_pointer == 111 && y_pointer == 85)
||(x_pointer == 112 && y_pointer == 85)
||(x_pointer == 113 && y_pointer == 85)
||(x_pointer == 114 && y_pointer == 85)
||(x_pointer == 115 && y_pointer == 85)
||(x_pointer == 116 && y_pointer == 85)
||(x_pointer == 117 && y_pointer == 85)
||(x_pointer == 118 && y_pointer == 85)
||(x_pointer == 5 && y_pointer == 86)
||(x_pointer == 6 && y_pointer == 86)
||(x_pointer == 7 && y_pointer == 86)
||(x_pointer == 8 && y_pointer == 86)
||(x_pointer == 9 && y_pointer == 86)
||(x_pointer == 10 && y_pointer == 86)
||(x_pointer == 11 && y_pointer == 86)
||(x_pointer == 12 && y_pointer == 86)
||(x_pointer == 13 && y_pointer == 86)
||(x_pointer == 14 && y_pointer == 86)
||(x_pointer == 15 && y_pointer == 86)
||(x_pointer == 16 && y_pointer == 86)
||(x_pointer == 17 && y_pointer == 86)
||(x_pointer == 18 && y_pointer == 86)
||(x_pointer == 19 && y_pointer == 86)
||(x_pointer == 20 && y_pointer == 86)
||(x_pointer == 21 && y_pointer == 86)
||(x_pointer == 22 && y_pointer == 86)
||(x_pointer == 23 && y_pointer == 86)
||(x_pointer == 24 && y_pointer == 86)
||(x_pointer == 25 && y_pointer == 86)
||(x_pointer == 26 && y_pointer == 86)
||(x_pointer == 27 && y_pointer == 86)
||(x_pointer == 28 && y_pointer == 86)
||(x_pointer == 29 && y_pointer == 86)
||(x_pointer == 30 && y_pointer == 86)
||(x_pointer == 31 && y_pointer == 86)
||(x_pointer == 32 && y_pointer == 86)
||(x_pointer == 33 && y_pointer == 86)
||(x_pointer == 34 && y_pointer == 86)
||(x_pointer == 35 && y_pointer == 86)
||(x_pointer == 36 && y_pointer == 86)
||(x_pointer == 37 && y_pointer == 86)
||(x_pointer == 38 && y_pointer == 86)
||(x_pointer == 39 && y_pointer == 86)
||(x_pointer == 40 && y_pointer == 86)
||(x_pointer == 41 && y_pointer == 86)
||(x_pointer == 42 && y_pointer == 86)
||(x_pointer == 43 && y_pointer == 86)
||(x_pointer == 44 && y_pointer == 86)
||(x_pointer == 45 && y_pointer == 86)
||(x_pointer == 46 && y_pointer == 86)
||(x_pointer == 47 && y_pointer == 86)
||(x_pointer == 48 && y_pointer == 86)
||(x_pointer == 49 && y_pointer == 86)
||(x_pointer == 50 && y_pointer == 86)
||(x_pointer == 51 && y_pointer == 86)
||(x_pointer == 52 && y_pointer == 86)
||(x_pointer == 53 && y_pointer == 86)
||(x_pointer == 54 && y_pointer == 86)
||(x_pointer == 55 && y_pointer == 86)
||(x_pointer == 56 && y_pointer == 86)
||(x_pointer == 57 && y_pointer == 86)
||(x_pointer == 58 && y_pointer == 86)
||(x_pointer == 110 && y_pointer == 86)
||(x_pointer == 111 && y_pointer == 86)
||(x_pointer == 112 && y_pointer == 86)
||(x_pointer == 113 && y_pointer == 86)
||(x_pointer == 114 && y_pointer == 86)
||(x_pointer == 115 && y_pointer == 86)
||(x_pointer == 116 && y_pointer == 86)
||(x_pointer == 117 && y_pointer == 86)
||(x_pointer == 118 && y_pointer == 86)
||(x_pointer == 5 && y_pointer == 87)
||(x_pointer == 6 && y_pointer == 87)
||(x_pointer == 7 && y_pointer == 87)
||(x_pointer == 8 && y_pointer == 87)
||(x_pointer == 9 && y_pointer == 87)
||(x_pointer == 10 && y_pointer == 87)
||(x_pointer == 11 && y_pointer == 87)
||(x_pointer == 12 && y_pointer == 87)
||(x_pointer == 13 && y_pointer == 87)
||(x_pointer == 14 && y_pointer == 87)
||(x_pointer == 15 && y_pointer == 87)
||(x_pointer == 16 && y_pointer == 87)
||(x_pointer == 17 && y_pointer == 87)
||(x_pointer == 18 && y_pointer == 87)
||(x_pointer == 19 && y_pointer == 87)
||(x_pointer == 20 && y_pointer == 87)
||(x_pointer == 21 && y_pointer == 87)
||(x_pointer == 22 && y_pointer == 87)
||(x_pointer == 23 && y_pointer == 87)
||(x_pointer == 24 && y_pointer == 87)
||(x_pointer == 25 && y_pointer == 87)
||(x_pointer == 26 && y_pointer == 87)
||(x_pointer == 27 && y_pointer == 87)
||(x_pointer == 28 && y_pointer == 87)
||(x_pointer == 29 && y_pointer == 87)
||(x_pointer == 30 && y_pointer == 87)
||(x_pointer == 31 && y_pointer == 87)
||(x_pointer == 32 && y_pointer == 87)
||(x_pointer == 33 && y_pointer == 87)
||(x_pointer == 34 && y_pointer == 87)
||(x_pointer == 35 && y_pointer == 87)
||(x_pointer == 36 && y_pointer == 87)
||(x_pointer == 37 && y_pointer == 87)
||(x_pointer == 38 && y_pointer == 87)
||(x_pointer == 39 && y_pointer == 87)
||(x_pointer == 40 && y_pointer == 87)
||(x_pointer == 41 && y_pointer == 87)
||(x_pointer == 42 && y_pointer == 87)
||(x_pointer == 43 && y_pointer == 87)
||(x_pointer == 44 && y_pointer == 87)
||(x_pointer == 45 && y_pointer == 87)
||(x_pointer == 46 && y_pointer == 87)
||(x_pointer == 47 && y_pointer == 87)
||(x_pointer == 48 && y_pointer == 87)
||(x_pointer == 49 && y_pointer == 87)
||(x_pointer == 50 && y_pointer == 87)
||(x_pointer == 51 && y_pointer == 87)
||(x_pointer == 52 && y_pointer == 87)
||(x_pointer == 53 && y_pointer == 87)
||(x_pointer == 54 && y_pointer == 87)
||(x_pointer == 55 && y_pointer == 87)
||(x_pointer == 56 && y_pointer == 87)
||(x_pointer == 57 && y_pointer == 87)
||(x_pointer == 58 && y_pointer == 87)
||(x_pointer == 110 && y_pointer == 87)
||(x_pointer == 111 && y_pointer == 87)
||(x_pointer == 112 && y_pointer == 87)
||(x_pointer == 113 && y_pointer == 87)
||(x_pointer == 114 && y_pointer == 87)
||(x_pointer == 115 && y_pointer == 87)
||(x_pointer == 116 && y_pointer == 87)
||(x_pointer == 117 && y_pointer == 87)
||(x_pointer == 118 && y_pointer == 87)
||(x_pointer == 5 && y_pointer == 88)
||(x_pointer == 6 && y_pointer == 88)
||(x_pointer == 7 && y_pointer == 88)
||(x_pointer == 8 && y_pointer == 88)
||(x_pointer == 9 && y_pointer == 88)
||(x_pointer == 10 && y_pointer == 88)
||(x_pointer == 11 && y_pointer == 88)
||(x_pointer == 12 && y_pointer == 88)
||(x_pointer == 13 && y_pointer == 88)
||(x_pointer == 14 && y_pointer == 88)
||(x_pointer == 15 && y_pointer == 88)
||(x_pointer == 16 && y_pointer == 88)
||(x_pointer == 17 && y_pointer == 88)
||(x_pointer == 18 && y_pointer == 88)
||(x_pointer == 19 && y_pointer == 88)
||(x_pointer == 20 && y_pointer == 88)
||(x_pointer == 21 && y_pointer == 88)
||(x_pointer == 22 && y_pointer == 88)
||(x_pointer == 23 && y_pointer == 88)
||(x_pointer == 24 && y_pointer == 88)
||(x_pointer == 25 && y_pointer == 88)
||(x_pointer == 26 && y_pointer == 88)
||(x_pointer == 27 && y_pointer == 88)
||(x_pointer == 28 && y_pointer == 88)
||(x_pointer == 29 && y_pointer == 88)
||(x_pointer == 30 && y_pointer == 88)
||(x_pointer == 31 && y_pointer == 88)
||(x_pointer == 32 && y_pointer == 88)
||(x_pointer == 33 && y_pointer == 88)
||(x_pointer == 34 && y_pointer == 88)
||(x_pointer == 35 && y_pointer == 88)
||(x_pointer == 36 && y_pointer == 88)
||(x_pointer == 37 && y_pointer == 88)
||(x_pointer == 38 && y_pointer == 88)
||(x_pointer == 39 && y_pointer == 88)
||(x_pointer == 40 && y_pointer == 88)
||(x_pointer == 41 && y_pointer == 88)
||(x_pointer == 42 && y_pointer == 88)
||(x_pointer == 43 && y_pointer == 88)
||(x_pointer == 44 && y_pointer == 88)
||(x_pointer == 45 && y_pointer == 88)
||(x_pointer == 46 && y_pointer == 88)
||(x_pointer == 47 && y_pointer == 88)
||(x_pointer == 48 && y_pointer == 88)
||(x_pointer == 49 && y_pointer == 88)
||(x_pointer == 50 && y_pointer == 88)
||(x_pointer == 51 && y_pointer == 88)
||(x_pointer == 52 && y_pointer == 88)
||(x_pointer == 53 && y_pointer == 88)
||(x_pointer == 54 && y_pointer == 88)
||(x_pointer == 55 && y_pointer == 88)
||(x_pointer == 56 && y_pointer == 88)
||(x_pointer == 57 && y_pointer == 88)
||(x_pointer == 58 && y_pointer == 88)
||(x_pointer == 110 && y_pointer == 88)
||(x_pointer == 111 && y_pointer == 88)
||(x_pointer == 112 && y_pointer == 88)
||(x_pointer == 113 && y_pointer == 88)
||(x_pointer == 114 && y_pointer == 88)
||(x_pointer == 115 && y_pointer == 88)
||(x_pointer == 116 && y_pointer == 88)
||(x_pointer == 117 && y_pointer == 88)
||(x_pointer == 118 && y_pointer == 88)
||(x_pointer == 5 && y_pointer == 89)
||(x_pointer == 6 && y_pointer == 89)
||(x_pointer == 7 && y_pointer == 89)
||(x_pointer == 8 && y_pointer == 89)
||(x_pointer == 9 && y_pointer == 89)
||(x_pointer == 10 && y_pointer == 89)
||(x_pointer == 11 && y_pointer == 89)
||(x_pointer == 12 && y_pointer == 89)
||(x_pointer == 13 && y_pointer == 89)
||(x_pointer == 14 && y_pointer == 89)
||(x_pointer == 15 && y_pointer == 89)
||(x_pointer == 16 && y_pointer == 89)
||(x_pointer == 17 && y_pointer == 89)
||(x_pointer == 18 && y_pointer == 89)
||(x_pointer == 19 && y_pointer == 89)
||(x_pointer == 20 && y_pointer == 89)
||(x_pointer == 21 && y_pointer == 89)
||(x_pointer == 22 && y_pointer == 89)
||(x_pointer == 23 && y_pointer == 89)
||(x_pointer == 24 && y_pointer == 89)
||(x_pointer == 25 && y_pointer == 89)
||(x_pointer == 26 && y_pointer == 89)
||(x_pointer == 27 && y_pointer == 89)
||(x_pointer == 28 && y_pointer == 89)
||(x_pointer == 29 && y_pointer == 89)
||(x_pointer == 30 && y_pointer == 89)
||(x_pointer == 31 && y_pointer == 89)
||(x_pointer == 32 && y_pointer == 89)
||(x_pointer == 33 && y_pointer == 89)
||(x_pointer == 34 && y_pointer == 89)
||(x_pointer == 35 && y_pointer == 89)
||(x_pointer == 36 && y_pointer == 89)
||(x_pointer == 37 && y_pointer == 89)
||(x_pointer == 38 && y_pointer == 89)
||(x_pointer == 39 && y_pointer == 89)
||(x_pointer == 40 && y_pointer == 89)
||(x_pointer == 41 && y_pointer == 89)
||(x_pointer == 42 && y_pointer == 89)
||(x_pointer == 43 && y_pointer == 89)
||(x_pointer == 44 && y_pointer == 89)
||(x_pointer == 45 && y_pointer == 89)
||(x_pointer == 46 && y_pointer == 89)
||(x_pointer == 47 && y_pointer == 89)
||(x_pointer == 48 && y_pointer == 89)
||(x_pointer == 49 && y_pointer == 89)
||(x_pointer == 50 && y_pointer == 89)
||(x_pointer == 51 && y_pointer == 89)
||(x_pointer == 52 && y_pointer == 89)
||(x_pointer == 53 && y_pointer == 89)
||(x_pointer == 54 && y_pointer == 89)
||(x_pointer == 55 && y_pointer == 89)
||(x_pointer == 56 && y_pointer == 89)
||(x_pointer == 57 && y_pointer == 89)
||(x_pointer == 58 && y_pointer == 89)
||(x_pointer == 110 && y_pointer == 89)
||(x_pointer == 111 && y_pointer == 89)
||(x_pointer == 112 && y_pointer == 89)
||(x_pointer == 113 && y_pointer == 89)
||(x_pointer == 114 && y_pointer == 89)
||(x_pointer == 115 && y_pointer == 89)
||(x_pointer == 116 && y_pointer == 89)
||(x_pointer == 117 && y_pointer == 89)
||(x_pointer == 118 && y_pointer == 89)
||(x_pointer == 5 && y_pointer == 90)
||(x_pointer == 6 && y_pointer == 90)
||(x_pointer == 7 && y_pointer == 90)
||(x_pointer == 8 && y_pointer == 90)
||(x_pointer == 9 && y_pointer == 90)
||(x_pointer == 10 && y_pointer == 90)
||(x_pointer == 11 && y_pointer == 90)
||(x_pointer == 12 && y_pointer == 90)
||(x_pointer == 13 && y_pointer == 90)
||(x_pointer == 14 && y_pointer == 90)
||(x_pointer == 15 && y_pointer == 90)
||(x_pointer == 16 && y_pointer == 90)
||(x_pointer == 17 && y_pointer == 90)
||(x_pointer == 18 && y_pointer == 90)
||(x_pointer == 19 && y_pointer == 90)
||(x_pointer == 20 && y_pointer == 90)
||(x_pointer == 21 && y_pointer == 90)
||(x_pointer == 22 && y_pointer == 90)
||(x_pointer == 23 && y_pointer == 90)
||(x_pointer == 24 && y_pointer == 90)
||(x_pointer == 25 && y_pointer == 90)
||(x_pointer == 26 && y_pointer == 90)
||(x_pointer == 27 && y_pointer == 90)
||(x_pointer == 28 && y_pointer == 90)
||(x_pointer == 29 && y_pointer == 90)
||(x_pointer == 30 && y_pointer == 90)
||(x_pointer == 31 && y_pointer == 90)
||(x_pointer == 32 && y_pointer == 90)
||(x_pointer == 33 && y_pointer == 90)
||(x_pointer == 34 && y_pointer == 90)
||(x_pointer == 35 && y_pointer == 90)
||(x_pointer == 36 && y_pointer == 90)
||(x_pointer == 37 && y_pointer == 90)
||(x_pointer == 38 && y_pointer == 90)
||(x_pointer == 39 && y_pointer == 90)
||(x_pointer == 40 && y_pointer == 90)
||(x_pointer == 41 && y_pointer == 90)
||(x_pointer == 42 && y_pointer == 90)
||(x_pointer == 43 && y_pointer == 90)
||(x_pointer == 44 && y_pointer == 90)
||(x_pointer == 45 && y_pointer == 90)
||(x_pointer == 46 && y_pointer == 90)
||(x_pointer == 47 && y_pointer == 90)
||(x_pointer == 48 && y_pointer == 90)
||(x_pointer == 49 && y_pointer == 90)
||(x_pointer == 50 && y_pointer == 90)
||(x_pointer == 51 && y_pointer == 90)
||(x_pointer == 52 && y_pointer == 90)
||(x_pointer == 53 && y_pointer == 90)
||(x_pointer == 54 && y_pointer == 90)
||(x_pointer == 55 && y_pointer == 90)
||(x_pointer == 56 && y_pointer == 90)
||(x_pointer == 57 && y_pointer == 90)
||(x_pointer == 58 && y_pointer == 90)
||(x_pointer == 110 && y_pointer == 90)
||(x_pointer == 111 && y_pointer == 90)
||(x_pointer == 112 && y_pointer == 90)
||(x_pointer == 113 && y_pointer == 90)
||(x_pointer == 114 && y_pointer == 90)
||(x_pointer == 115 && y_pointer == 90)
||(x_pointer == 116 && y_pointer == 90)
||(x_pointer == 117 && y_pointer == 90)
||(x_pointer == 118 && y_pointer == 90)
||(x_pointer == 5 && y_pointer == 91)
||(x_pointer == 6 && y_pointer == 91)
||(x_pointer == 7 && y_pointer == 91)
||(x_pointer == 8 && y_pointer == 91)
||(x_pointer == 9 && y_pointer == 91)
||(x_pointer == 10 && y_pointer == 91)
||(x_pointer == 11 && y_pointer == 91)
||(x_pointer == 12 && y_pointer == 91)
||(x_pointer == 13 && y_pointer == 91)
||(x_pointer == 14 && y_pointer == 91)
||(x_pointer == 15 && y_pointer == 91)
||(x_pointer == 16 && y_pointer == 91)
||(x_pointer == 17 && y_pointer == 91)
||(x_pointer == 18 && y_pointer == 91)
||(x_pointer == 19 && y_pointer == 91)
||(x_pointer == 20 && y_pointer == 91)
||(x_pointer == 21 && y_pointer == 91)
||(x_pointer == 22 && y_pointer == 91)
||(x_pointer == 23 && y_pointer == 91)
||(x_pointer == 24 && y_pointer == 91)
||(x_pointer == 25 && y_pointer == 91)
||(x_pointer == 26 && y_pointer == 91)
||(x_pointer == 27 && y_pointer == 91)
||(x_pointer == 28 && y_pointer == 91)
||(x_pointer == 29 && y_pointer == 91)
||(x_pointer == 30 && y_pointer == 91)
||(x_pointer == 31 && y_pointer == 91)
||(x_pointer == 32 && y_pointer == 91)
||(x_pointer == 33 && y_pointer == 91)
||(x_pointer == 34 && y_pointer == 91)
||(x_pointer == 35 && y_pointer == 91)
||(x_pointer == 36 && y_pointer == 91)
||(x_pointer == 37 && y_pointer == 91)
||(x_pointer == 38 && y_pointer == 91)
||(x_pointer == 39 && y_pointer == 91)
||(x_pointer == 40 && y_pointer == 91)
||(x_pointer == 41 && y_pointer == 91)
||(x_pointer == 42 && y_pointer == 91)
||(x_pointer == 43 && y_pointer == 91)
||(x_pointer == 44 && y_pointer == 91)
||(x_pointer == 45 && y_pointer == 91)
||(x_pointer == 46 && y_pointer == 91)
||(x_pointer == 47 && y_pointer == 91)
||(x_pointer == 48 && y_pointer == 91)
||(x_pointer == 49 && y_pointer == 91)
||(x_pointer == 50 && y_pointer == 91)
||(x_pointer == 51 && y_pointer == 91)
||(x_pointer == 52 && y_pointer == 91)
||(x_pointer == 53 && y_pointer == 91)
||(x_pointer == 54 && y_pointer == 91)
||(x_pointer == 55 && y_pointer == 91)
||(x_pointer == 56 && y_pointer == 91)
||(x_pointer == 57 && y_pointer == 91)
||(x_pointer == 58 && y_pointer == 91)
||(x_pointer == 110 && y_pointer == 91)
||(x_pointer == 111 && y_pointer == 91)
||(x_pointer == 112 && y_pointer == 91)
||(x_pointer == 113 && y_pointer == 91)
||(x_pointer == 114 && y_pointer == 91)
||(x_pointer == 115 && y_pointer == 91)
||(x_pointer == 116 && y_pointer == 91)
||(x_pointer == 117 && y_pointer == 91)
||(x_pointer == 118 && y_pointer == 91)
||(x_pointer == 5 && y_pointer == 92)
||(x_pointer == 6 && y_pointer == 92)
||(x_pointer == 7 && y_pointer == 92)
||(x_pointer == 8 && y_pointer == 92)
||(x_pointer == 9 && y_pointer == 92)
||(x_pointer == 10 && y_pointer == 92)
||(x_pointer == 11 && y_pointer == 92)
||(x_pointer == 12 && y_pointer == 92)
||(x_pointer == 13 && y_pointer == 92)
||(x_pointer == 14 && y_pointer == 92)
||(x_pointer == 15 && y_pointer == 92)
||(x_pointer == 16 && y_pointer == 92)
||(x_pointer == 17 && y_pointer == 92)
||(x_pointer == 18 && y_pointer == 92)
||(x_pointer == 19 && y_pointer == 92)
||(x_pointer == 20 && y_pointer == 92)
||(x_pointer == 21 && y_pointer == 92)
||(x_pointer == 22 && y_pointer == 92)
||(x_pointer == 23 && y_pointer == 92)
||(x_pointer == 24 && y_pointer == 92)
||(x_pointer == 25 && y_pointer == 92)
||(x_pointer == 26 && y_pointer == 92)
||(x_pointer == 27 && y_pointer == 92)
||(x_pointer == 28 && y_pointer == 92)
||(x_pointer == 29 && y_pointer == 92)
||(x_pointer == 30 && y_pointer == 92)
||(x_pointer == 31 && y_pointer == 92)
||(x_pointer == 32 && y_pointer == 92)
||(x_pointer == 33 && y_pointer == 92)
||(x_pointer == 34 && y_pointer == 92)
||(x_pointer == 35 && y_pointer == 92)
||(x_pointer == 36 && y_pointer == 92)
||(x_pointer == 37 && y_pointer == 92)
||(x_pointer == 38 && y_pointer == 92)
||(x_pointer == 39 && y_pointer == 92)
||(x_pointer == 40 && y_pointer == 92)
||(x_pointer == 41 && y_pointer == 92)
||(x_pointer == 42 && y_pointer == 92)
||(x_pointer == 43 && y_pointer == 92)
||(x_pointer == 44 && y_pointer == 92)
||(x_pointer == 45 && y_pointer == 92)
||(x_pointer == 46 && y_pointer == 92)
||(x_pointer == 47 && y_pointer == 92)
||(x_pointer == 48 && y_pointer == 92)
||(x_pointer == 49 && y_pointer == 92)
||(x_pointer == 50 && y_pointer == 92)
||(x_pointer == 51 && y_pointer == 92)
||(x_pointer == 52 && y_pointer == 92)
||(x_pointer == 53 && y_pointer == 92)
||(x_pointer == 54 && y_pointer == 92)
||(x_pointer == 55 && y_pointer == 92)
||(x_pointer == 56 && y_pointer == 92)
||(x_pointer == 57 && y_pointer == 92)
||(x_pointer == 58 && y_pointer == 92)
||(x_pointer == 110 && y_pointer == 92)
||(x_pointer == 111 && y_pointer == 92)
||(x_pointer == 112 && y_pointer == 92)
||(x_pointer == 113 && y_pointer == 92)
||(x_pointer == 114 && y_pointer == 92)
||(x_pointer == 115 && y_pointer == 92)
||(x_pointer == 116 && y_pointer == 92)
||(x_pointer == 117 && y_pointer == 92)
||(x_pointer == 118 && y_pointer == 92)
||(x_pointer == 5 && y_pointer == 93)
||(x_pointer == 6 && y_pointer == 93)
||(x_pointer == 7 && y_pointer == 93)
||(x_pointer == 8 && y_pointer == 93)
||(x_pointer == 9 && y_pointer == 93)
||(x_pointer == 10 && y_pointer == 93)
||(x_pointer == 11 && y_pointer == 93)
||(x_pointer == 12 && y_pointer == 93)
||(x_pointer == 13 && y_pointer == 93)
||(x_pointer == 14 && y_pointer == 93)
||(x_pointer == 15 && y_pointer == 93)
||(x_pointer == 16 && y_pointer == 93)
||(x_pointer == 17 && y_pointer == 93)
||(x_pointer == 18 && y_pointer == 93)
||(x_pointer == 19 && y_pointer == 93)
||(x_pointer == 20 && y_pointer == 93)
||(x_pointer == 21 && y_pointer == 93)
||(x_pointer == 22 && y_pointer == 93)
||(x_pointer == 23 && y_pointer == 93)
||(x_pointer == 24 && y_pointer == 93)
||(x_pointer == 25 && y_pointer == 93)
||(x_pointer == 26 && y_pointer == 93)
||(x_pointer == 27 && y_pointer == 93)
||(x_pointer == 28 && y_pointer == 93)
||(x_pointer == 29 && y_pointer == 93)
||(x_pointer == 30 && y_pointer == 93)
||(x_pointer == 31 && y_pointer == 93)
||(x_pointer == 32 && y_pointer == 93)
||(x_pointer == 33 && y_pointer == 93)
||(x_pointer == 34 && y_pointer == 93)
||(x_pointer == 35 && y_pointer == 93)
||(x_pointer == 36 && y_pointer == 93)
||(x_pointer == 37 && y_pointer == 93)
||(x_pointer == 38 && y_pointer == 93)
||(x_pointer == 39 && y_pointer == 93)
||(x_pointer == 40 && y_pointer == 93)
||(x_pointer == 41 && y_pointer == 93)
||(x_pointer == 42 && y_pointer == 93)
||(x_pointer == 43 && y_pointer == 93)
||(x_pointer == 44 && y_pointer == 93)
||(x_pointer == 45 && y_pointer == 93)
||(x_pointer == 46 && y_pointer == 93)
||(x_pointer == 47 && y_pointer == 93)
||(x_pointer == 48 && y_pointer == 93)
||(x_pointer == 49 && y_pointer == 93)
||(x_pointer == 50 && y_pointer == 93)
||(x_pointer == 51 && y_pointer == 93)
||(x_pointer == 52 && y_pointer == 93)
||(x_pointer == 53 && y_pointer == 93)
||(x_pointer == 54 && y_pointer == 93)
||(x_pointer == 55 && y_pointer == 93)
||(x_pointer == 56 && y_pointer == 93)
||(x_pointer == 57 && y_pointer == 93)
||(x_pointer == 58 && y_pointer == 93)
||(x_pointer == 110 && y_pointer == 93)
||(x_pointer == 111 && y_pointer == 93)
||(x_pointer == 112 && y_pointer == 93)
||(x_pointer == 113 && y_pointer == 93)
||(x_pointer == 114 && y_pointer == 93)
||(x_pointer == 115 && y_pointer == 93)
||(x_pointer == 116 && y_pointer == 93)
||(x_pointer == 117 && y_pointer == 93)
||(x_pointer == 118 && y_pointer == 93)
||(x_pointer == 5 && y_pointer == 94)
||(x_pointer == 6 && y_pointer == 94)
||(x_pointer == 7 && y_pointer == 94)
||(x_pointer == 8 && y_pointer == 94)
||(x_pointer == 9 && y_pointer == 94)
||(x_pointer == 10 && y_pointer == 94)
||(x_pointer == 11 && y_pointer == 94)
||(x_pointer == 12 && y_pointer == 94)
||(x_pointer == 13 && y_pointer == 94)
||(x_pointer == 14 && y_pointer == 94)
||(x_pointer == 15 && y_pointer == 94)
||(x_pointer == 16 && y_pointer == 94)
||(x_pointer == 17 && y_pointer == 94)
||(x_pointer == 18 && y_pointer == 94)
||(x_pointer == 19 && y_pointer == 94)
||(x_pointer == 20 && y_pointer == 94)
||(x_pointer == 21 && y_pointer == 94)
||(x_pointer == 22 && y_pointer == 94)
||(x_pointer == 23 && y_pointer == 94)
||(x_pointer == 24 && y_pointer == 94)
||(x_pointer == 25 && y_pointer == 94)
||(x_pointer == 26 && y_pointer == 94)
||(x_pointer == 27 && y_pointer == 94)
||(x_pointer == 28 && y_pointer == 94)
||(x_pointer == 29 && y_pointer == 94)
||(x_pointer == 30 && y_pointer == 94)
||(x_pointer == 31 && y_pointer == 94)
||(x_pointer == 32 && y_pointer == 94)
||(x_pointer == 33 && y_pointer == 94)
||(x_pointer == 34 && y_pointer == 94)
||(x_pointer == 35 && y_pointer == 94)
||(x_pointer == 36 && y_pointer == 94)
||(x_pointer == 37 && y_pointer == 94)
||(x_pointer == 38 && y_pointer == 94)
||(x_pointer == 39 && y_pointer == 94)
||(x_pointer == 40 && y_pointer == 94)
||(x_pointer == 41 && y_pointer == 94)
||(x_pointer == 42 && y_pointer == 94)
||(x_pointer == 43 && y_pointer == 94)
||(x_pointer == 44 && y_pointer == 94)
||(x_pointer == 45 && y_pointer == 94)
||(x_pointer == 46 && y_pointer == 94)
||(x_pointer == 47 && y_pointer == 94)
||(x_pointer == 48 && y_pointer == 94)
||(x_pointer == 49 && y_pointer == 94)
||(x_pointer == 50 && y_pointer == 94)
||(x_pointer == 51 && y_pointer == 94)
||(x_pointer == 52 && y_pointer == 94)
||(x_pointer == 53 && y_pointer == 94)
||(x_pointer == 54 && y_pointer == 94)
||(x_pointer == 55 && y_pointer == 94)
||(x_pointer == 56 && y_pointer == 94)
||(x_pointer == 57 && y_pointer == 94)
||(x_pointer == 58 && y_pointer == 94)
||(x_pointer == 110 && y_pointer == 94)
||(x_pointer == 111 && y_pointer == 94)
||(x_pointer == 112 && y_pointer == 94)
||(x_pointer == 113 && y_pointer == 94)
||(x_pointer == 114 && y_pointer == 94)
||(x_pointer == 115 && y_pointer == 94)
||(x_pointer == 116 && y_pointer == 94)
||(x_pointer == 117 && y_pointer == 94)
||(x_pointer == 118 && y_pointer == 94)
||(x_pointer == 110 && y_pointer == 95)
||(x_pointer == 111 && y_pointer == 95)
||(x_pointer == 112 && y_pointer == 95)
||(x_pointer == 113 && y_pointer == 95)
||(x_pointer == 114 && y_pointer == 95)
||(x_pointer == 115 && y_pointer == 95)
||(x_pointer == 116 && y_pointer == 95)
||(x_pointer == 117 && y_pointer == 95)
||(x_pointer == 118 && y_pointer == 95)
||(x_pointer == 110 && y_pointer == 96)
||(x_pointer == 111 && y_pointer == 96)
||(x_pointer == 112 && y_pointer == 96)
||(x_pointer == 113 && y_pointer == 96)
||(x_pointer == 114 && y_pointer == 96)
||(x_pointer == 115 && y_pointer == 96)
||(x_pointer == 116 && y_pointer == 96)
||(x_pointer == 117 && y_pointer == 96)
||(x_pointer == 118 && y_pointer == 96)
||(x_pointer == 110 && y_pointer == 97)
||(x_pointer == 111 && y_pointer == 97)
||(x_pointer == 112 && y_pointer == 97)
||(x_pointer == 113 && y_pointer == 97)
||(x_pointer == 114 && y_pointer == 97)
||(x_pointer == 115 && y_pointer == 97)
||(x_pointer == 116 && y_pointer == 97)
||(x_pointer == 117 && y_pointer == 97)
||(x_pointer == 118 && y_pointer == 97)
||(x_pointer == 110 && y_pointer == 98)
||(x_pointer == 111 && y_pointer == 98)
||(x_pointer == 112 && y_pointer == 98)
||(x_pointer == 113 && y_pointer == 98)
||(x_pointer == 114 && y_pointer == 98)
||(x_pointer == 115 && y_pointer == 98)
||(x_pointer == 116 && y_pointer == 98)
||(x_pointer == 117 && y_pointer == 98)
||(x_pointer == 118 && y_pointer == 98)
||(x_pointer == 110 && y_pointer == 99)
||(x_pointer == 111 && y_pointer == 99)
||(x_pointer == 112 && y_pointer == 99)
||(x_pointer == 113 && y_pointer == 99)
||(x_pointer == 114 && y_pointer == 99)
||(x_pointer == 115 && y_pointer == 99)
||(x_pointer == 116 && y_pointer == 99)
||(x_pointer == 117 && y_pointer == 99)
||(x_pointer == 118 && y_pointer == 99)
||(x_pointer == 110 && y_pointer == 100)
||(x_pointer == 111 && y_pointer == 100)
||(x_pointer == 112 && y_pointer == 100)
||(x_pointer == 113 && y_pointer == 100)
||(x_pointer == 114 && y_pointer == 100)
||(x_pointer == 115 && y_pointer == 100)
||(x_pointer == 116 && y_pointer == 100)
||(x_pointer == 117 && y_pointer == 100)
||(x_pointer == 118 && y_pointer == 100)
||(x_pointer == 110 && y_pointer == 101)
||(x_pointer == 111 && y_pointer == 101)
||(x_pointer == 112 && y_pointer == 101)
||(x_pointer == 113 && y_pointer == 101)
||(x_pointer == 114 && y_pointer == 101)
||(x_pointer == 115 && y_pointer == 101)
||(x_pointer == 116 && y_pointer == 101)
||(x_pointer == 117 && y_pointer == 101)
||(x_pointer == 118 && y_pointer == 101)
||(x_pointer == 110 && y_pointer == 102)
||(x_pointer == 111 && y_pointer == 102)
||(x_pointer == 112 && y_pointer == 102)
||(x_pointer == 113 && y_pointer == 102)
||(x_pointer == 114 && y_pointer == 102)
||(x_pointer == 115 && y_pointer == 102)
||(x_pointer == 116 && y_pointer == 102)
||(x_pointer == 117 && y_pointer == 102)
||(x_pointer == 118 && y_pointer == 102)
||(x_pointer == 110 && y_pointer == 103)
||(x_pointer == 111 && y_pointer == 103)
||(x_pointer == 112 && y_pointer == 103)
||(x_pointer == 113 && y_pointer == 103)
||(x_pointer == 114 && y_pointer == 103)
||(x_pointer == 115 && y_pointer == 103)
||(x_pointer == 116 && y_pointer == 103)
||(x_pointer == 117 && y_pointer == 103)
||(x_pointer == 118 && y_pointer == 103)
||(x_pointer == 71 && y_pointer == 104)
||(x_pointer == 72 && y_pointer == 104)
||(x_pointer == 73 && y_pointer == 104)
||(x_pointer == 74 && y_pointer == 104)
||(x_pointer == 75 && y_pointer == 104)
||(x_pointer == 76 && y_pointer == 104)
||(x_pointer == 77 && y_pointer == 104)
||(x_pointer == 78 && y_pointer == 104)
||(x_pointer == 79 && y_pointer == 104)
||(x_pointer == 80 && y_pointer == 104)
||(x_pointer == 81 && y_pointer == 104)
||(x_pointer == 82 && y_pointer == 104)
||(x_pointer == 83 && y_pointer == 104)
||(x_pointer == 84 && y_pointer == 104)
||(x_pointer == 85 && y_pointer == 104)
||(x_pointer == 86 && y_pointer == 104)
||(x_pointer == 87 && y_pointer == 104)
||(x_pointer == 88 && y_pointer == 104)
||(x_pointer == 89 && y_pointer == 104)
||(x_pointer == 90 && y_pointer == 104)
||(x_pointer == 91 && y_pointer == 104)
||(x_pointer == 92 && y_pointer == 104)
||(x_pointer == 93 && y_pointer == 104)
||(x_pointer == 94 && y_pointer == 104)
||(x_pointer == 95 && y_pointer == 104)
||(x_pointer == 96 && y_pointer == 104)
||(x_pointer == 97 && y_pointer == 104)
||(x_pointer == 98 && y_pointer == 104)
||(x_pointer == 99 && y_pointer == 104)
||(x_pointer == 100 && y_pointer == 104)
||(x_pointer == 101 && y_pointer == 104)
||(x_pointer == 102 && y_pointer == 104)
||(x_pointer == 103 && y_pointer == 104)
||(x_pointer == 104 && y_pointer == 104)
||(x_pointer == 105 && y_pointer == 104)
||(x_pointer == 106 && y_pointer == 104)
||(x_pointer == 107 && y_pointer == 104)
||(x_pointer == 108 && y_pointer == 104)
||(x_pointer == 109 && y_pointer == 104)
||(x_pointer == 110 && y_pointer == 104)
||(x_pointer == 111 && y_pointer == 104)
||(x_pointer == 112 && y_pointer == 104)
||(x_pointer == 113 && y_pointer == 104)
||(x_pointer == 114 && y_pointer == 104)
||(x_pointer == 115 && y_pointer == 104)
||(x_pointer == 116 && y_pointer == 104)
||(x_pointer == 117 && y_pointer == 104)
||(x_pointer == 118 && y_pointer == 104)
||(x_pointer == 119 && y_pointer == 104)
||(x_pointer == 120 && y_pointer == 104)
||(x_pointer == 121 && y_pointer == 104)
||(x_pointer == 122 && y_pointer == 104)
||(x_pointer == 123 && y_pointer == 104)
||(x_pointer == 124 && y_pointer == 104)
||(x_pointer == 125 && y_pointer == 104)
||(x_pointer == 126 && y_pointer == 104)
||(x_pointer == 127 && y_pointer == 104)
||(x_pointer == 128 && y_pointer == 104)
||(x_pointer == 129 && y_pointer == 104)
||(x_pointer == 130 && y_pointer == 104)
||(x_pointer == 131 && y_pointer == 104)
||(x_pointer == 132 && y_pointer == 104)
||(x_pointer == 133 && y_pointer == 104)
||(x_pointer == 134 && y_pointer == 104)
||(x_pointer == 135 && y_pointer == 104)
||(x_pointer == 136 && y_pointer == 104)
||(x_pointer == 137 && y_pointer == 104)
||(x_pointer == 138 && y_pointer == 104)
||(x_pointer == 139 && y_pointer == 104)
||(x_pointer == 140 && y_pointer == 104)
||(x_pointer == 141 && y_pointer == 104)
||(x_pointer == 142 && y_pointer == 104)
||(x_pointer == 143 && y_pointer == 104)
||(x_pointer == 144 && y_pointer == 104)
||(x_pointer == 145 && y_pointer == 104)
||(x_pointer == 146 && y_pointer == 104)
||(x_pointer == 147 && y_pointer == 104)
||(x_pointer == 148 && y_pointer == 104)
||(x_pointer == 149 && y_pointer == 104)
||(x_pointer == 150 && y_pointer == 104)
||(x_pointer == 151 && y_pointer == 104)
||(x_pointer == 152 && y_pointer == 104)
||(x_pointer == 153 && y_pointer == 104)
||(x_pointer == 154 && y_pointer == 104)
||(x_pointer == 71 && y_pointer == 105)
||(x_pointer == 72 && y_pointer == 105)
||(x_pointer == 73 && y_pointer == 105)
||(x_pointer == 74 && y_pointer == 105)
||(x_pointer == 75 && y_pointer == 105)
||(x_pointer == 76 && y_pointer == 105)
||(x_pointer == 77 && y_pointer == 105)
||(x_pointer == 78 && y_pointer == 105)
||(x_pointer == 79 && y_pointer == 105)
||(x_pointer == 80 && y_pointer == 105)
||(x_pointer == 81 && y_pointer == 105)
||(x_pointer == 82 && y_pointer == 105)
||(x_pointer == 83 && y_pointer == 105)
||(x_pointer == 84 && y_pointer == 105)
||(x_pointer == 85 && y_pointer == 105)
||(x_pointer == 86 && y_pointer == 105)
||(x_pointer == 87 && y_pointer == 105)
||(x_pointer == 88 && y_pointer == 105)
||(x_pointer == 89 && y_pointer == 105)
||(x_pointer == 90 && y_pointer == 105)
||(x_pointer == 91 && y_pointer == 105)
||(x_pointer == 92 && y_pointer == 105)
||(x_pointer == 93 && y_pointer == 105)
||(x_pointer == 94 && y_pointer == 105)
||(x_pointer == 95 && y_pointer == 105)
||(x_pointer == 96 && y_pointer == 105)
||(x_pointer == 97 && y_pointer == 105)
||(x_pointer == 98 && y_pointer == 105)
||(x_pointer == 99 && y_pointer == 105)
||(x_pointer == 100 && y_pointer == 105)
||(x_pointer == 101 && y_pointer == 105)
||(x_pointer == 102 && y_pointer == 105)
||(x_pointer == 103 && y_pointer == 105)
||(x_pointer == 104 && y_pointer == 105)
||(x_pointer == 105 && y_pointer == 105)
||(x_pointer == 106 && y_pointer == 105)
||(x_pointer == 107 && y_pointer == 105)
||(x_pointer == 108 && y_pointer == 105)
||(x_pointer == 109 && y_pointer == 105)
||(x_pointer == 110 && y_pointer == 105)
||(x_pointer == 111 && y_pointer == 105)
||(x_pointer == 112 && y_pointer == 105)
||(x_pointer == 113 && y_pointer == 105)
||(x_pointer == 114 && y_pointer == 105)
||(x_pointer == 115 && y_pointer == 105)
||(x_pointer == 116 && y_pointer == 105)
||(x_pointer == 117 && y_pointer == 105)
||(x_pointer == 118 && y_pointer == 105)
||(x_pointer == 119 && y_pointer == 105)
||(x_pointer == 120 && y_pointer == 105)
||(x_pointer == 121 && y_pointer == 105)
||(x_pointer == 122 && y_pointer == 105)
||(x_pointer == 123 && y_pointer == 105)
||(x_pointer == 124 && y_pointer == 105)
||(x_pointer == 125 && y_pointer == 105)
||(x_pointer == 126 && y_pointer == 105)
||(x_pointer == 127 && y_pointer == 105)
||(x_pointer == 128 && y_pointer == 105)
||(x_pointer == 129 && y_pointer == 105)
||(x_pointer == 130 && y_pointer == 105)
||(x_pointer == 131 && y_pointer == 105)
||(x_pointer == 132 && y_pointer == 105)
||(x_pointer == 133 && y_pointer == 105)
||(x_pointer == 134 && y_pointer == 105)
||(x_pointer == 135 && y_pointer == 105)
||(x_pointer == 136 && y_pointer == 105)
||(x_pointer == 137 && y_pointer == 105)
||(x_pointer == 138 && y_pointer == 105)
||(x_pointer == 139 && y_pointer == 105)
||(x_pointer == 140 && y_pointer == 105)
||(x_pointer == 141 && y_pointer == 105)
||(x_pointer == 142 && y_pointer == 105)
||(x_pointer == 143 && y_pointer == 105)
||(x_pointer == 144 && y_pointer == 105)
||(x_pointer == 145 && y_pointer == 105)
||(x_pointer == 146 && y_pointer == 105)
||(x_pointer == 147 && y_pointer == 105)
||(x_pointer == 148 && y_pointer == 105)
||(x_pointer == 149 && y_pointer == 105)
||(x_pointer == 150 && y_pointer == 105)
||(x_pointer == 151 && y_pointer == 105)
||(x_pointer == 152 && y_pointer == 105)
||(x_pointer == 153 && y_pointer == 105)
||(x_pointer == 154 && y_pointer == 105)
||(x_pointer == 71 && y_pointer == 106)
||(x_pointer == 72 && y_pointer == 106)
||(x_pointer == 73 && y_pointer == 106)
||(x_pointer == 74 && y_pointer == 106)
||(x_pointer == 75 && y_pointer == 106)
||(x_pointer == 76 && y_pointer == 106)
||(x_pointer == 77 && y_pointer == 106)
||(x_pointer == 78 && y_pointer == 106)
||(x_pointer == 79 && y_pointer == 106)
||(x_pointer == 80 && y_pointer == 106)
||(x_pointer == 81 && y_pointer == 106)
||(x_pointer == 82 && y_pointer == 106)
||(x_pointer == 83 && y_pointer == 106)
||(x_pointer == 84 && y_pointer == 106)
||(x_pointer == 85 && y_pointer == 106)
||(x_pointer == 86 && y_pointer == 106)
||(x_pointer == 87 && y_pointer == 106)
||(x_pointer == 88 && y_pointer == 106)
||(x_pointer == 89 && y_pointer == 106)
||(x_pointer == 90 && y_pointer == 106)
||(x_pointer == 91 && y_pointer == 106)
||(x_pointer == 92 && y_pointer == 106)
||(x_pointer == 93 && y_pointer == 106)
||(x_pointer == 94 && y_pointer == 106)
||(x_pointer == 95 && y_pointer == 106)
||(x_pointer == 96 && y_pointer == 106)
||(x_pointer == 97 && y_pointer == 106)
||(x_pointer == 98 && y_pointer == 106)
||(x_pointer == 99 && y_pointer == 106)
||(x_pointer == 100 && y_pointer == 106)
||(x_pointer == 101 && y_pointer == 106)
||(x_pointer == 102 && y_pointer == 106)
||(x_pointer == 103 && y_pointer == 106)
||(x_pointer == 104 && y_pointer == 106)
||(x_pointer == 105 && y_pointer == 106)
||(x_pointer == 106 && y_pointer == 106)
||(x_pointer == 107 && y_pointer == 106)
||(x_pointer == 108 && y_pointer == 106)
||(x_pointer == 109 && y_pointer == 106)
||(x_pointer == 110 && y_pointer == 106)
||(x_pointer == 111 && y_pointer == 106)
||(x_pointer == 112 && y_pointer == 106)
||(x_pointer == 113 && y_pointer == 106)
||(x_pointer == 114 && y_pointer == 106)
||(x_pointer == 115 && y_pointer == 106)
||(x_pointer == 116 && y_pointer == 106)
||(x_pointer == 117 && y_pointer == 106)
||(x_pointer == 118 && y_pointer == 106)
||(x_pointer == 119 && y_pointer == 106)
||(x_pointer == 120 && y_pointer == 106)
||(x_pointer == 121 && y_pointer == 106)
||(x_pointer == 122 && y_pointer == 106)
||(x_pointer == 123 && y_pointer == 106)
||(x_pointer == 124 && y_pointer == 106)
||(x_pointer == 125 && y_pointer == 106)
||(x_pointer == 126 && y_pointer == 106)
||(x_pointer == 127 && y_pointer == 106)
||(x_pointer == 128 && y_pointer == 106)
||(x_pointer == 129 && y_pointer == 106)
||(x_pointer == 130 && y_pointer == 106)
||(x_pointer == 131 && y_pointer == 106)
||(x_pointer == 132 && y_pointer == 106)
||(x_pointer == 133 && y_pointer == 106)
||(x_pointer == 134 && y_pointer == 106)
||(x_pointer == 135 && y_pointer == 106)
||(x_pointer == 136 && y_pointer == 106)
||(x_pointer == 137 && y_pointer == 106)
||(x_pointer == 138 && y_pointer == 106)
||(x_pointer == 139 && y_pointer == 106)
||(x_pointer == 140 && y_pointer == 106)
||(x_pointer == 141 && y_pointer == 106)
||(x_pointer == 142 && y_pointer == 106)
||(x_pointer == 143 && y_pointer == 106)
||(x_pointer == 144 && y_pointer == 106)
||(x_pointer == 145 && y_pointer == 106)
||(x_pointer == 146 && y_pointer == 106)
||(x_pointer == 147 && y_pointer == 106)
||(x_pointer == 148 && y_pointer == 106)
||(x_pointer == 149 && y_pointer == 106)
||(x_pointer == 150 && y_pointer == 106)
||(x_pointer == 151 && y_pointer == 106)
||(x_pointer == 152 && y_pointer == 106)
||(x_pointer == 153 && y_pointer == 106)
||(x_pointer == 154 && y_pointer == 106)
||(x_pointer == 71 && y_pointer == 107)
||(x_pointer == 72 && y_pointer == 107)
||(x_pointer == 73 && y_pointer == 107)
||(x_pointer == 74 && y_pointer == 107)
||(x_pointer == 75 && y_pointer == 107)
||(x_pointer == 76 && y_pointer == 107)
||(x_pointer == 77 && y_pointer == 107)
||(x_pointer == 78 && y_pointer == 107)
||(x_pointer == 79 && y_pointer == 107)
||(x_pointer == 80 && y_pointer == 107)
||(x_pointer == 81 && y_pointer == 107)
||(x_pointer == 82 && y_pointer == 107)
||(x_pointer == 83 && y_pointer == 107)
||(x_pointer == 84 && y_pointer == 107)
||(x_pointer == 85 && y_pointer == 107)
||(x_pointer == 86 && y_pointer == 107)
||(x_pointer == 87 && y_pointer == 107)
||(x_pointer == 88 && y_pointer == 107)
||(x_pointer == 89 && y_pointer == 107)
||(x_pointer == 90 && y_pointer == 107)
||(x_pointer == 91 && y_pointer == 107)
||(x_pointer == 92 && y_pointer == 107)
||(x_pointer == 93 && y_pointer == 107)
||(x_pointer == 94 && y_pointer == 107)
||(x_pointer == 95 && y_pointer == 107)
||(x_pointer == 96 && y_pointer == 107)
||(x_pointer == 97 && y_pointer == 107)
||(x_pointer == 98 && y_pointer == 107)
||(x_pointer == 99 && y_pointer == 107)
||(x_pointer == 100 && y_pointer == 107)
||(x_pointer == 101 && y_pointer == 107)
||(x_pointer == 102 && y_pointer == 107)
||(x_pointer == 103 && y_pointer == 107)
||(x_pointer == 104 && y_pointer == 107)
||(x_pointer == 105 && y_pointer == 107)
||(x_pointer == 106 && y_pointer == 107)
||(x_pointer == 107 && y_pointer == 107)
||(x_pointer == 108 && y_pointer == 107)
||(x_pointer == 109 && y_pointer == 107)
||(x_pointer == 110 && y_pointer == 107)
||(x_pointer == 111 && y_pointer == 107)
||(x_pointer == 112 && y_pointer == 107)
||(x_pointer == 113 && y_pointer == 107)
||(x_pointer == 114 && y_pointer == 107)
||(x_pointer == 115 && y_pointer == 107)
||(x_pointer == 116 && y_pointer == 107)
||(x_pointer == 117 && y_pointer == 107)
||(x_pointer == 118 && y_pointer == 107)
||(x_pointer == 119 && y_pointer == 107)
||(x_pointer == 120 && y_pointer == 107)
||(x_pointer == 121 && y_pointer == 107)
||(x_pointer == 122 && y_pointer == 107)
||(x_pointer == 123 && y_pointer == 107)
||(x_pointer == 124 && y_pointer == 107)
||(x_pointer == 125 && y_pointer == 107)
||(x_pointer == 126 && y_pointer == 107)
||(x_pointer == 127 && y_pointer == 107)
||(x_pointer == 128 && y_pointer == 107)
||(x_pointer == 129 && y_pointer == 107)
||(x_pointer == 130 && y_pointer == 107)
||(x_pointer == 131 && y_pointer == 107)
||(x_pointer == 132 && y_pointer == 107)
||(x_pointer == 133 && y_pointer == 107)
||(x_pointer == 134 && y_pointer == 107)
||(x_pointer == 135 && y_pointer == 107)
||(x_pointer == 136 && y_pointer == 107)
||(x_pointer == 137 && y_pointer == 107)
||(x_pointer == 138 && y_pointer == 107)
||(x_pointer == 139 && y_pointer == 107)
||(x_pointer == 140 && y_pointer == 107)
||(x_pointer == 141 && y_pointer == 107)
||(x_pointer == 142 && y_pointer == 107)
||(x_pointer == 143 && y_pointer == 107)
||(x_pointer == 144 && y_pointer == 107)
||(x_pointer == 145 && y_pointer == 107)
||(x_pointer == 146 && y_pointer == 107)
||(x_pointer == 147 && y_pointer == 107)
||(x_pointer == 148 && y_pointer == 107)
||(x_pointer == 149 && y_pointer == 107)
||(x_pointer == 150 && y_pointer == 107)
||(x_pointer == 151 && y_pointer == 107)
||(x_pointer == 152 && y_pointer == 107)
||(x_pointer == 153 && y_pointer == 107)
||(x_pointer == 154 && y_pointer == 107)
||(x_pointer == 71 && y_pointer == 108)
||(x_pointer == 72 && y_pointer == 108)
||(x_pointer == 73 && y_pointer == 108)
||(x_pointer == 74 && y_pointer == 108)
||(x_pointer == 75 && y_pointer == 108)
||(x_pointer == 76 && y_pointer == 108)
||(x_pointer == 77 && y_pointer == 108)
||(x_pointer == 78 && y_pointer == 108)
||(x_pointer == 79 && y_pointer == 108)
||(x_pointer == 80 && y_pointer == 108)
||(x_pointer == 81 && y_pointer == 108)
||(x_pointer == 82 && y_pointer == 108)
||(x_pointer == 83 && y_pointer == 108)
||(x_pointer == 84 && y_pointer == 108)
||(x_pointer == 85 && y_pointer == 108)
||(x_pointer == 86 && y_pointer == 108)
||(x_pointer == 87 && y_pointer == 108)
||(x_pointer == 88 && y_pointer == 108)
||(x_pointer == 89 && y_pointer == 108)
||(x_pointer == 90 && y_pointer == 108)
||(x_pointer == 91 && y_pointer == 108)
||(x_pointer == 92 && y_pointer == 108)
||(x_pointer == 93 && y_pointer == 108)
||(x_pointer == 94 && y_pointer == 108)
||(x_pointer == 95 && y_pointer == 108)
||(x_pointer == 96 && y_pointer == 108)
||(x_pointer == 97 && y_pointer == 108)
||(x_pointer == 98 && y_pointer == 108)
||(x_pointer == 99 && y_pointer == 108)
||(x_pointer == 100 && y_pointer == 108)
||(x_pointer == 101 && y_pointer == 108)
||(x_pointer == 102 && y_pointer == 108)
||(x_pointer == 103 && y_pointer == 108)
||(x_pointer == 104 && y_pointer == 108)
||(x_pointer == 105 && y_pointer == 108)
||(x_pointer == 106 && y_pointer == 108)
||(x_pointer == 107 && y_pointer == 108)
||(x_pointer == 108 && y_pointer == 108)
||(x_pointer == 109 && y_pointer == 108)
||(x_pointer == 110 && y_pointer == 108)
||(x_pointer == 111 && y_pointer == 108)
||(x_pointer == 112 && y_pointer == 108)
||(x_pointer == 113 && y_pointer == 108)
||(x_pointer == 114 && y_pointer == 108)
||(x_pointer == 115 && y_pointer == 108)
||(x_pointer == 116 && y_pointer == 108)
||(x_pointer == 117 && y_pointer == 108)
||(x_pointer == 118 && y_pointer == 108)
||(x_pointer == 119 && y_pointer == 108)
||(x_pointer == 120 && y_pointer == 108)
||(x_pointer == 121 && y_pointer == 108)
||(x_pointer == 122 && y_pointer == 108)
||(x_pointer == 123 && y_pointer == 108)
||(x_pointer == 124 && y_pointer == 108)
||(x_pointer == 125 && y_pointer == 108)
||(x_pointer == 126 && y_pointer == 108)
||(x_pointer == 127 && y_pointer == 108)
||(x_pointer == 128 && y_pointer == 108)
||(x_pointer == 129 && y_pointer == 108)
||(x_pointer == 130 && y_pointer == 108)
||(x_pointer == 131 && y_pointer == 108)
||(x_pointer == 132 && y_pointer == 108)
||(x_pointer == 133 && y_pointer == 108)
||(x_pointer == 134 && y_pointer == 108)
||(x_pointer == 135 && y_pointer == 108)
||(x_pointer == 136 && y_pointer == 108)
||(x_pointer == 137 && y_pointer == 108)
||(x_pointer == 138 && y_pointer == 108)
||(x_pointer == 139 && y_pointer == 108)
||(x_pointer == 140 && y_pointer == 108)
||(x_pointer == 141 && y_pointer == 108)
||(x_pointer == 142 && y_pointer == 108)
||(x_pointer == 143 && y_pointer == 108)
||(x_pointer == 144 && y_pointer == 108)
||(x_pointer == 145 && y_pointer == 108)
||(x_pointer == 146 && y_pointer == 108)
||(x_pointer == 147 && y_pointer == 108)
||(x_pointer == 148 && y_pointer == 108)
||(x_pointer == 149 && y_pointer == 108)
||(x_pointer == 150 && y_pointer == 108)
||(x_pointer == 151 && y_pointer == 108)
||(x_pointer == 152 && y_pointer == 108)
||(x_pointer == 153 && y_pointer == 108)
||(x_pointer == 154 && y_pointer == 108)
||(x_pointer == 71 && y_pointer == 109)
||(x_pointer == 72 && y_pointer == 109)
||(x_pointer == 73 && y_pointer == 109)
||(x_pointer == 74 && y_pointer == 109)
||(x_pointer == 75 && y_pointer == 109)
||(x_pointer == 76 && y_pointer == 109)
||(x_pointer == 77 && y_pointer == 109)
||(x_pointer == 78 && y_pointer == 109)
||(x_pointer == 79 && y_pointer == 109)
||(x_pointer == 80 && y_pointer == 109)
||(x_pointer == 81 && y_pointer == 109)
||(x_pointer == 82 && y_pointer == 109)
||(x_pointer == 83 && y_pointer == 109)
||(x_pointer == 84 && y_pointer == 109)
||(x_pointer == 85 && y_pointer == 109)
||(x_pointer == 86 && y_pointer == 109)
||(x_pointer == 87 && y_pointer == 109)
||(x_pointer == 88 && y_pointer == 109)
||(x_pointer == 89 && y_pointer == 109)
||(x_pointer == 90 && y_pointer == 109)
||(x_pointer == 91 && y_pointer == 109)
||(x_pointer == 92 && y_pointer == 109)
||(x_pointer == 93 && y_pointer == 109)
||(x_pointer == 94 && y_pointer == 109)
||(x_pointer == 95 && y_pointer == 109)
||(x_pointer == 96 && y_pointer == 109)
||(x_pointer == 97 && y_pointer == 109)
||(x_pointer == 98 && y_pointer == 109)
||(x_pointer == 99 && y_pointer == 109)
||(x_pointer == 100 && y_pointer == 109)
||(x_pointer == 101 && y_pointer == 109)
||(x_pointer == 102 && y_pointer == 109)
||(x_pointer == 103 && y_pointer == 109)
||(x_pointer == 104 && y_pointer == 109)
||(x_pointer == 105 && y_pointer == 109)
||(x_pointer == 106 && y_pointer == 109)
||(x_pointer == 107 && y_pointer == 109)
||(x_pointer == 108 && y_pointer == 109)
||(x_pointer == 109 && y_pointer == 109)
||(x_pointer == 110 && y_pointer == 109)
||(x_pointer == 111 && y_pointer == 109)
||(x_pointer == 112 && y_pointer == 109)
||(x_pointer == 113 && y_pointer == 109)
||(x_pointer == 114 && y_pointer == 109)
||(x_pointer == 115 && y_pointer == 109)
||(x_pointer == 116 && y_pointer == 109)
||(x_pointer == 117 && y_pointer == 109)
||(x_pointer == 118 && y_pointer == 109)
||(x_pointer == 119 && y_pointer == 109)
||(x_pointer == 120 && y_pointer == 109)
||(x_pointer == 121 && y_pointer == 109)
||(x_pointer == 122 && y_pointer == 109)
||(x_pointer == 123 && y_pointer == 109)
||(x_pointer == 124 && y_pointer == 109)
||(x_pointer == 125 && y_pointer == 109)
||(x_pointer == 126 && y_pointer == 109)
||(x_pointer == 127 && y_pointer == 109)
||(x_pointer == 128 && y_pointer == 109)
||(x_pointer == 129 && y_pointer == 109)
||(x_pointer == 130 && y_pointer == 109)
||(x_pointer == 131 && y_pointer == 109)
||(x_pointer == 132 && y_pointer == 109)
||(x_pointer == 133 && y_pointer == 109)
||(x_pointer == 134 && y_pointer == 109)
||(x_pointer == 135 && y_pointer == 109)
||(x_pointer == 136 && y_pointer == 109)
||(x_pointer == 137 && y_pointer == 109)
||(x_pointer == 138 && y_pointer == 109)
||(x_pointer == 139 && y_pointer == 109)
||(x_pointer == 140 && y_pointer == 109)
||(x_pointer == 141 && y_pointer == 109)
||(x_pointer == 142 && y_pointer == 109)
||(x_pointer == 143 && y_pointer == 109)
||(x_pointer == 144 && y_pointer == 109)
||(x_pointer == 145 && y_pointer == 109)
||(x_pointer == 146 && y_pointer == 109)
||(x_pointer == 147 && y_pointer == 109)
||(x_pointer == 148 && y_pointer == 109)
||(x_pointer == 149 && y_pointer == 109)
||(x_pointer == 150 && y_pointer == 109)
||(x_pointer == 151 && y_pointer == 109)
||(x_pointer == 152 && y_pointer == 109)
||(x_pointer == 153 && y_pointer == 109)
||(x_pointer == 154 && y_pointer == 109));
	
	
	wire barrier_pixel_5 = current_level == 5 && ((x_pointer == 2 && y_pointer == 2)
||(x_pointer == 3 && y_pointer == 2)
||(x_pointer == 4 && y_pointer == 2)
||(x_pointer == 5 && y_pointer == 2)
||(x_pointer == 6 && y_pointer == 2)
||(x_pointer == 7 && y_pointer == 2)
||(x_pointer == 8 && y_pointer == 2)
||(x_pointer == 9 && y_pointer == 2)
||(x_pointer == 10 && y_pointer == 2)
||(x_pointer == 11 && y_pointer == 2)
||(x_pointer == 12 && y_pointer == 2)
||(x_pointer == 13 && y_pointer == 2)
||(x_pointer == 14 && y_pointer == 2)
||(x_pointer == 15 && y_pointer == 2)
||(x_pointer == 16 && y_pointer == 2)
||(x_pointer == 17 && y_pointer == 2)
||(x_pointer == 18 && y_pointer == 2)
||(x_pointer == 19 && y_pointer == 2)
||(x_pointer == 20 && y_pointer == 2)
||(x_pointer == 21 && y_pointer == 2)
||(x_pointer == 22 && y_pointer == 2)
||(x_pointer == 23 && y_pointer == 2)
||(x_pointer == 24 && y_pointer == 2)
||(x_pointer == 25 && y_pointer == 2)
||(x_pointer == 26 && y_pointer == 2)
||(x_pointer == 27 && y_pointer == 2)
||(x_pointer == 28 && y_pointer == 2)
||(x_pointer == 29 && y_pointer == 2)
||(x_pointer == 30 && y_pointer == 2)
||(x_pointer == 31 && y_pointer == 2)
||(x_pointer == 32 && y_pointer == 2)
||(x_pointer == 33 && y_pointer == 2)
||(x_pointer == 34 && y_pointer == 2)
||(x_pointer == 35 && y_pointer == 2)
||(x_pointer == 36 && y_pointer == 2)
||(x_pointer == 37 && y_pointer == 2)
||(x_pointer == 38 && y_pointer == 2)
||(x_pointer == 39 && y_pointer == 2)
||(x_pointer == 40 && y_pointer == 2)
||(x_pointer == 41 && y_pointer == 2)
||(x_pointer == 42 && y_pointer == 2)
||(x_pointer == 43 && y_pointer == 2)
||(x_pointer == 44 && y_pointer == 2)
||(x_pointer == 45 && y_pointer == 2)
||(x_pointer == 46 && y_pointer == 2)
||(x_pointer == 47 && y_pointer == 2)
||(x_pointer == 48 && y_pointer == 2)
||(x_pointer == 49 && y_pointer == 2)
||(x_pointer == 50 && y_pointer == 2)
||(x_pointer == 51 && y_pointer == 2)
||(x_pointer == 52 && y_pointer == 2)
||(x_pointer == 53 && y_pointer == 2)
||(x_pointer == 54 && y_pointer == 2)
||(x_pointer == 55 && y_pointer == 2)
||(x_pointer == 56 && y_pointer == 2)
||(x_pointer == 57 && y_pointer == 2)
||(x_pointer == 58 && y_pointer == 2)
||(x_pointer == 59 && y_pointer == 2)
||(x_pointer == 60 && y_pointer == 2)
||(x_pointer == 61 && y_pointer == 2)
||(x_pointer == 62 && y_pointer == 2)
||(x_pointer == 63 && y_pointer == 2)
||(x_pointer == 64 && y_pointer == 2)
||(x_pointer == 65 && y_pointer == 2)
||(x_pointer == 66 && y_pointer == 2)
||(x_pointer == 67 && y_pointer == 2)
||(x_pointer == 68 && y_pointer == 2)
||(x_pointer == 69 && y_pointer == 2)
||(x_pointer == 70 && y_pointer == 2)
||(x_pointer == 71 && y_pointer == 2)
||(x_pointer == 72 && y_pointer == 2)
||(x_pointer == 73 && y_pointer == 2)
||(x_pointer == 74 && y_pointer == 2)
||(x_pointer == 75 && y_pointer == 2)
||(x_pointer == 76 && y_pointer == 2)
||(x_pointer == 77 && y_pointer == 2)
||(x_pointer == 78 && y_pointer == 2)
||(x_pointer == 79 && y_pointer == 2)
||(x_pointer == 80 && y_pointer == 2)
||(x_pointer == 81 && y_pointer == 2)
||(x_pointer == 82 && y_pointer == 2)
||(x_pointer == 83 && y_pointer == 2)
||(x_pointer == 84 && y_pointer == 2)
||(x_pointer == 85 && y_pointer == 2)
||(x_pointer == 86 && y_pointer == 2)
||(x_pointer == 87 && y_pointer == 2)
||(x_pointer == 88 && y_pointer == 2)
||(x_pointer == 89 && y_pointer == 2)
||(x_pointer == 90 && y_pointer == 2)
||(x_pointer == 91 && y_pointer == 2)
||(x_pointer == 92 && y_pointer == 2)
||(x_pointer == 93 && y_pointer == 2)
||(x_pointer == 94 && y_pointer == 2)
||(x_pointer == 95 && y_pointer == 2)
||(x_pointer == 96 && y_pointer == 2)
||(x_pointer == 97 && y_pointer == 2)
||(x_pointer == 98 && y_pointer == 2)
||(x_pointer == 99 && y_pointer == 2)
||(x_pointer == 100 && y_pointer == 2)
||(x_pointer == 101 && y_pointer == 2)
||(x_pointer == 102 && y_pointer == 2)
||(x_pointer == 103 && y_pointer == 2)
||(x_pointer == 104 && y_pointer == 2)
||(x_pointer == 105 && y_pointer == 2)
||(x_pointer == 106 && y_pointer == 2)
||(x_pointer == 107 && y_pointer == 2)
||(x_pointer == 108 && y_pointer == 2)
||(x_pointer == 109 && y_pointer == 2)
||(x_pointer == 110 && y_pointer == 2)
||(x_pointer == 111 && y_pointer == 2)
||(x_pointer == 112 && y_pointer == 2)
||(x_pointer == 113 && y_pointer == 2)
||(x_pointer == 114 && y_pointer == 2)
||(x_pointer == 115 && y_pointer == 2)
||(x_pointer == 116 && y_pointer == 2)
||(x_pointer == 117 && y_pointer == 2)
||(x_pointer == 118 && y_pointer == 2)
||(x_pointer == 119 && y_pointer == 2)
||(x_pointer == 120 && y_pointer == 2)
||(x_pointer == 121 && y_pointer == 2)
||(x_pointer == 122 && y_pointer == 2)
||(x_pointer == 123 && y_pointer == 2)
||(x_pointer == 124 && y_pointer == 2)
||(x_pointer == 125 && y_pointer == 2)
||(x_pointer == 126 && y_pointer == 2)
||(x_pointer == 127 && y_pointer == 2)
||(x_pointer == 128 && y_pointer == 2)
||(x_pointer == 129 && y_pointer == 2)
||(x_pointer == 130 && y_pointer == 2)
||(x_pointer == 131 && y_pointer == 2)
||(x_pointer == 132 && y_pointer == 2)
||(x_pointer == 133 && y_pointer == 2)
||(x_pointer == 134 && y_pointer == 2)
||(x_pointer == 135 && y_pointer == 2)
||(x_pointer == 136 && y_pointer == 2)
||(x_pointer == 137 && y_pointer == 2)
||(x_pointer == 138 && y_pointer == 2)
||(x_pointer == 139 && y_pointer == 2)
||(x_pointer == 140 && y_pointer == 2)
||(x_pointer == 141 && y_pointer == 2)
||(x_pointer == 142 && y_pointer == 2)
||(x_pointer == 143 && y_pointer == 2)
||(x_pointer == 144 && y_pointer == 2)
||(x_pointer == 145 && y_pointer == 2)
||(x_pointer == 146 && y_pointer == 2)
||(x_pointer == 147 && y_pointer == 2)
||(x_pointer == 148 && y_pointer == 2)
||(x_pointer == 149 && y_pointer == 2)
||(x_pointer == 150 && y_pointer == 2)
||(x_pointer == 151 && y_pointer == 2)
||(x_pointer == 152 && y_pointer == 2)
||(x_pointer == 153 && y_pointer == 2)
||(x_pointer == 154 && y_pointer == 2)
||(x_pointer == 155 && y_pointer == 2)
||(x_pointer == 156 && y_pointer == 2)
||(x_pointer == 157 && y_pointer == 2)
||(x_pointer == 2 && y_pointer == 3)
||(x_pointer == 3 && y_pointer == 3)
||(x_pointer == 4 && y_pointer == 3)
||(x_pointer == 5 && y_pointer == 3)
||(x_pointer == 6 && y_pointer == 3)
||(x_pointer == 7 && y_pointer == 3)
||(x_pointer == 8 && y_pointer == 3)
||(x_pointer == 9 && y_pointer == 3)
||(x_pointer == 10 && y_pointer == 3)
||(x_pointer == 11 && y_pointer == 3)
||(x_pointer == 12 && y_pointer == 3)
||(x_pointer == 13 && y_pointer == 3)
||(x_pointer == 14 && y_pointer == 3)
||(x_pointer == 15 && y_pointer == 3)
||(x_pointer == 16 && y_pointer == 3)
||(x_pointer == 17 && y_pointer == 3)
||(x_pointer == 18 && y_pointer == 3)
||(x_pointer == 19 && y_pointer == 3)
||(x_pointer == 20 && y_pointer == 3)
||(x_pointer == 21 && y_pointer == 3)
||(x_pointer == 22 && y_pointer == 3)
||(x_pointer == 23 && y_pointer == 3)
||(x_pointer == 24 && y_pointer == 3)
||(x_pointer == 25 && y_pointer == 3)
||(x_pointer == 26 && y_pointer == 3)
||(x_pointer == 27 && y_pointer == 3)
||(x_pointer == 28 && y_pointer == 3)
||(x_pointer == 29 && y_pointer == 3)
||(x_pointer == 30 && y_pointer == 3)
||(x_pointer == 31 && y_pointer == 3)
||(x_pointer == 32 && y_pointer == 3)
||(x_pointer == 33 && y_pointer == 3)
||(x_pointer == 34 && y_pointer == 3)
||(x_pointer == 35 && y_pointer == 3)
||(x_pointer == 36 && y_pointer == 3)
||(x_pointer == 37 && y_pointer == 3)
||(x_pointer == 38 && y_pointer == 3)
||(x_pointer == 39 && y_pointer == 3)
||(x_pointer == 40 && y_pointer == 3)
||(x_pointer == 41 && y_pointer == 3)
||(x_pointer == 42 && y_pointer == 3)
||(x_pointer == 43 && y_pointer == 3)
||(x_pointer == 44 && y_pointer == 3)
||(x_pointer == 45 && y_pointer == 3)
||(x_pointer == 46 && y_pointer == 3)
||(x_pointer == 47 && y_pointer == 3)
||(x_pointer == 48 && y_pointer == 3)
||(x_pointer == 49 && y_pointer == 3)
||(x_pointer == 50 && y_pointer == 3)
||(x_pointer == 51 && y_pointer == 3)
||(x_pointer == 52 && y_pointer == 3)
||(x_pointer == 53 && y_pointer == 3)
||(x_pointer == 54 && y_pointer == 3)
||(x_pointer == 55 && y_pointer == 3)
||(x_pointer == 56 && y_pointer == 3)
||(x_pointer == 57 && y_pointer == 3)
||(x_pointer == 58 && y_pointer == 3)
||(x_pointer == 59 && y_pointer == 3)
||(x_pointer == 60 && y_pointer == 3)
||(x_pointer == 61 && y_pointer == 3)
||(x_pointer == 62 && y_pointer == 3)
||(x_pointer == 63 && y_pointer == 3)
||(x_pointer == 64 && y_pointer == 3)
||(x_pointer == 65 && y_pointer == 3)
||(x_pointer == 66 && y_pointer == 3)
||(x_pointer == 67 && y_pointer == 3)
||(x_pointer == 68 && y_pointer == 3)
||(x_pointer == 69 && y_pointer == 3)
||(x_pointer == 70 && y_pointer == 3)
||(x_pointer == 71 && y_pointer == 3)
||(x_pointer == 72 && y_pointer == 3)
||(x_pointer == 73 && y_pointer == 3)
||(x_pointer == 74 && y_pointer == 3)
||(x_pointer == 75 && y_pointer == 3)
||(x_pointer == 76 && y_pointer == 3)
||(x_pointer == 77 && y_pointer == 3)
||(x_pointer == 78 && y_pointer == 3)
||(x_pointer == 79 && y_pointer == 3)
||(x_pointer == 80 && y_pointer == 3)
||(x_pointer == 81 && y_pointer == 3)
||(x_pointer == 82 && y_pointer == 3)
||(x_pointer == 83 && y_pointer == 3)
||(x_pointer == 84 && y_pointer == 3)
||(x_pointer == 85 && y_pointer == 3)
||(x_pointer == 86 && y_pointer == 3)
||(x_pointer == 87 && y_pointer == 3)
||(x_pointer == 88 && y_pointer == 3)
||(x_pointer == 89 && y_pointer == 3)
||(x_pointer == 90 && y_pointer == 3)
||(x_pointer == 91 && y_pointer == 3)
||(x_pointer == 92 && y_pointer == 3)
||(x_pointer == 93 && y_pointer == 3)
||(x_pointer == 94 && y_pointer == 3)
||(x_pointer == 95 && y_pointer == 3)
||(x_pointer == 96 && y_pointer == 3)
||(x_pointer == 97 && y_pointer == 3)
||(x_pointer == 98 && y_pointer == 3)
||(x_pointer == 99 && y_pointer == 3)
||(x_pointer == 100 && y_pointer == 3)
||(x_pointer == 101 && y_pointer == 3)
||(x_pointer == 102 && y_pointer == 3)
||(x_pointer == 103 && y_pointer == 3)
||(x_pointer == 104 && y_pointer == 3)
||(x_pointer == 105 && y_pointer == 3)
||(x_pointer == 106 && y_pointer == 3)
||(x_pointer == 107 && y_pointer == 3)
||(x_pointer == 108 && y_pointer == 3)
||(x_pointer == 109 && y_pointer == 3)
||(x_pointer == 110 && y_pointer == 3)
||(x_pointer == 111 && y_pointer == 3)
||(x_pointer == 112 && y_pointer == 3)
||(x_pointer == 113 && y_pointer == 3)
||(x_pointer == 114 && y_pointer == 3)
||(x_pointer == 115 && y_pointer == 3)
||(x_pointer == 116 && y_pointer == 3)
||(x_pointer == 117 && y_pointer == 3)
||(x_pointer == 118 && y_pointer == 3)
||(x_pointer == 119 && y_pointer == 3)
||(x_pointer == 120 && y_pointer == 3)
||(x_pointer == 121 && y_pointer == 3)
||(x_pointer == 122 && y_pointer == 3)
||(x_pointer == 123 && y_pointer == 3)
||(x_pointer == 124 && y_pointer == 3)
||(x_pointer == 125 && y_pointer == 3)
||(x_pointer == 126 && y_pointer == 3)
||(x_pointer == 127 && y_pointer == 3)
||(x_pointer == 128 && y_pointer == 3)
||(x_pointer == 129 && y_pointer == 3)
||(x_pointer == 130 && y_pointer == 3)
||(x_pointer == 131 && y_pointer == 3)
||(x_pointer == 132 && y_pointer == 3)
||(x_pointer == 133 && y_pointer == 3)
||(x_pointer == 134 && y_pointer == 3)
||(x_pointer == 135 && y_pointer == 3)
||(x_pointer == 136 && y_pointer == 3)
||(x_pointer == 137 && y_pointer == 3)
||(x_pointer == 138 && y_pointer == 3)
||(x_pointer == 139 && y_pointer == 3)
||(x_pointer == 140 && y_pointer == 3)
||(x_pointer == 141 && y_pointer == 3)
||(x_pointer == 142 && y_pointer == 3)
||(x_pointer == 143 && y_pointer == 3)
||(x_pointer == 144 && y_pointer == 3)
||(x_pointer == 145 && y_pointer == 3)
||(x_pointer == 146 && y_pointer == 3)
||(x_pointer == 147 && y_pointer == 3)
||(x_pointer == 148 && y_pointer == 3)
||(x_pointer == 149 && y_pointer == 3)
||(x_pointer == 150 && y_pointer == 3)
||(x_pointer == 151 && y_pointer == 3)
||(x_pointer == 152 && y_pointer == 3)
||(x_pointer == 153 && y_pointer == 3)
||(x_pointer == 154 && y_pointer == 3)
||(x_pointer == 155 && y_pointer == 3)
||(x_pointer == 156 && y_pointer == 3)
||(x_pointer == 157 && y_pointer == 3)
||(x_pointer == 2 && y_pointer == 4)
||(x_pointer == 3 && y_pointer == 4)
||(x_pointer == 4 && y_pointer == 4)
||(x_pointer == 5 && y_pointer == 4)
||(x_pointer == 6 && y_pointer == 4)
||(x_pointer == 7 && y_pointer == 4)
||(x_pointer == 8 && y_pointer == 4)
||(x_pointer == 9 && y_pointer == 4)
||(x_pointer == 10 && y_pointer == 4)
||(x_pointer == 11 && y_pointer == 4)
||(x_pointer == 12 && y_pointer == 4)
||(x_pointer == 13 && y_pointer == 4)
||(x_pointer == 14 && y_pointer == 4)
||(x_pointer == 15 && y_pointer == 4)
||(x_pointer == 16 && y_pointer == 4)
||(x_pointer == 17 && y_pointer == 4)
||(x_pointer == 18 && y_pointer == 4)
||(x_pointer == 19 && y_pointer == 4)
||(x_pointer == 20 && y_pointer == 4)
||(x_pointer == 21 && y_pointer == 4)
||(x_pointer == 22 && y_pointer == 4)
||(x_pointer == 23 && y_pointer == 4)
||(x_pointer == 24 && y_pointer == 4)
||(x_pointer == 25 && y_pointer == 4)
||(x_pointer == 26 && y_pointer == 4)
||(x_pointer == 27 && y_pointer == 4)
||(x_pointer == 28 && y_pointer == 4)
||(x_pointer == 29 && y_pointer == 4)
||(x_pointer == 30 && y_pointer == 4)
||(x_pointer == 31 && y_pointer == 4)
||(x_pointer == 32 && y_pointer == 4)
||(x_pointer == 33 && y_pointer == 4)
||(x_pointer == 34 && y_pointer == 4)
||(x_pointer == 35 && y_pointer == 4)
||(x_pointer == 36 && y_pointer == 4)
||(x_pointer == 37 && y_pointer == 4)
||(x_pointer == 38 && y_pointer == 4)
||(x_pointer == 39 && y_pointer == 4)
||(x_pointer == 40 && y_pointer == 4)
||(x_pointer == 41 && y_pointer == 4)
||(x_pointer == 42 && y_pointer == 4)
||(x_pointer == 43 && y_pointer == 4)
||(x_pointer == 44 && y_pointer == 4)
||(x_pointer == 45 && y_pointer == 4)
||(x_pointer == 46 && y_pointer == 4)
||(x_pointer == 47 && y_pointer == 4)
||(x_pointer == 48 && y_pointer == 4)
||(x_pointer == 49 && y_pointer == 4)
||(x_pointer == 50 && y_pointer == 4)
||(x_pointer == 51 && y_pointer == 4)
||(x_pointer == 52 && y_pointer == 4)
||(x_pointer == 53 && y_pointer == 4)
||(x_pointer == 54 && y_pointer == 4)
||(x_pointer == 55 && y_pointer == 4)
||(x_pointer == 56 && y_pointer == 4)
||(x_pointer == 57 && y_pointer == 4)
||(x_pointer == 58 && y_pointer == 4)
||(x_pointer == 59 && y_pointer == 4)
||(x_pointer == 60 && y_pointer == 4)
||(x_pointer == 61 && y_pointer == 4)
||(x_pointer == 62 && y_pointer == 4)
||(x_pointer == 63 && y_pointer == 4)
||(x_pointer == 64 && y_pointer == 4)
||(x_pointer == 65 && y_pointer == 4)
||(x_pointer == 66 && y_pointer == 4)
||(x_pointer == 67 && y_pointer == 4)
||(x_pointer == 68 && y_pointer == 4)
||(x_pointer == 69 && y_pointer == 4)
||(x_pointer == 70 && y_pointer == 4)
||(x_pointer == 71 && y_pointer == 4)
||(x_pointer == 72 && y_pointer == 4)
||(x_pointer == 73 && y_pointer == 4)
||(x_pointer == 74 && y_pointer == 4)
||(x_pointer == 75 && y_pointer == 4)
||(x_pointer == 76 && y_pointer == 4)
||(x_pointer == 77 && y_pointer == 4)
||(x_pointer == 78 && y_pointer == 4)
||(x_pointer == 79 && y_pointer == 4)
||(x_pointer == 80 && y_pointer == 4)
||(x_pointer == 81 && y_pointer == 4)
||(x_pointer == 82 && y_pointer == 4)
||(x_pointer == 83 && y_pointer == 4)
||(x_pointer == 84 && y_pointer == 4)
||(x_pointer == 85 && y_pointer == 4)
||(x_pointer == 86 && y_pointer == 4)
||(x_pointer == 87 && y_pointer == 4)
||(x_pointer == 88 && y_pointer == 4)
||(x_pointer == 89 && y_pointer == 4)
||(x_pointer == 90 && y_pointer == 4)
||(x_pointer == 91 && y_pointer == 4)
||(x_pointer == 92 && y_pointer == 4)
||(x_pointer == 93 && y_pointer == 4)
||(x_pointer == 94 && y_pointer == 4)
||(x_pointer == 95 && y_pointer == 4)
||(x_pointer == 96 && y_pointer == 4)
||(x_pointer == 97 && y_pointer == 4)
||(x_pointer == 98 && y_pointer == 4)
||(x_pointer == 99 && y_pointer == 4)
||(x_pointer == 100 && y_pointer == 4)
||(x_pointer == 101 && y_pointer == 4)
||(x_pointer == 102 && y_pointer == 4)
||(x_pointer == 103 && y_pointer == 4)
||(x_pointer == 104 && y_pointer == 4)
||(x_pointer == 105 && y_pointer == 4)
||(x_pointer == 106 && y_pointer == 4)
||(x_pointer == 107 && y_pointer == 4)
||(x_pointer == 108 && y_pointer == 4)
||(x_pointer == 109 && y_pointer == 4)
||(x_pointer == 110 && y_pointer == 4)
||(x_pointer == 111 && y_pointer == 4)
||(x_pointer == 112 && y_pointer == 4)
||(x_pointer == 113 && y_pointer == 4)
||(x_pointer == 114 && y_pointer == 4)
||(x_pointer == 115 && y_pointer == 4)
||(x_pointer == 116 && y_pointer == 4)
||(x_pointer == 117 && y_pointer == 4)
||(x_pointer == 118 && y_pointer == 4)
||(x_pointer == 119 && y_pointer == 4)
||(x_pointer == 120 && y_pointer == 4)
||(x_pointer == 121 && y_pointer == 4)
||(x_pointer == 122 && y_pointer == 4)
||(x_pointer == 123 && y_pointer == 4)
||(x_pointer == 124 && y_pointer == 4)
||(x_pointer == 125 && y_pointer == 4)
||(x_pointer == 126 && y_pointer == 4)
||(x_pointer == 127 && y_pointer == 4)
||(x_pointer == 128 && y_pointer == 4)
||(x_pointer == 129 && y_pointer == 4)
||(x_pointer == 130 && y_pointer == 4)
||(x_pointer == 131 && y_pointer == 4)
||(x_pointer == 132 && y_pointer == 4)
||(x_pointer == 133 && y_pointer == 4)
||(x_pointer == 134 && y_pointer == 4)
||(x_pointer == 135 && y_pointer == 4)
||(x_pointer == 136 && y_pointer == 4)
||(x_pointer == 137 && y_pointer == 4)
||(x_pointer == 138 && y_pointer == 4)
||(x_pointer == 139 && y_pointer == 4)
||(x_pointer == 140 && y_pointer == 4)
||(x_pointer == 141 && y_pointer == 4)
||(x_pointer == 142 && y_pointer == 4)
||(x_pointer == 143 && y_pointer == 4)
||(x_pointer == 144 && y_pointer == 4)
||(x_pointer == 145 && y_pointer == 4)
||(x_pointer == 146 && y_pointer == 4)
||(x_pointer == 147 && y_pointer == 4)
||(x_pointer == 148 && y_pointer == 4)
||(x_pointer == 149 && y_pointer == 4)
||(x_pointer == 150 && y_pointer == 4)
||(x_pointer == 151 && y_pointer == 4)
||(x_pointer == 152 && y_pointer == 4)
||(x_pointer == 153 && y_pointer == 4)
||(x_pointer == 154 && y_pointer == 4)
||(x_pointer == 155 && y_pointer == 4)
||(x_pointer == 156 && y_pointer == 4)
||(x_pointer == 157 && y_pointer == 4)
||(x_pointer == 2 && y_pointer == 5)
||(x_pointer == 3 && y_pointer == 5)
||(x_pointer == 4 && y_pointer == 5)
||(x_pointer == 155 && y_pointer == 5)
||(x_pointer == 156 && y_pointer == 5)
||(x_pointer == 157 && y_pointer == 5)
||(x_pointer == 2 && y_pointer == 6)
||(x_pointer == 3 && y_pointer == 6)
||(x_pointer == 4 && y_pointer == 6)
||(x_pointer == 155 && y_pointer == 6)
||(x_pointer == 156 && y_pointer == 6)
||(x_pointer == 157 && y_pointer == 6)
||(x_pointer == 2 && y_pointer == 7)
||(x_pointer == 3 && y_pointer == 7)
||(x_pointer == 4 && y_pointer == 7)
||(x_pointer == 155 && y_pointer == 7)
||(x_pointer == 156 && y_pointer == 7)
||(x_pointer == 157 && y_pointer == 7)
||(x_pointer == 2 && y_pointer == 8)
||(x_pointer == 3 && y_pointer == 8)
||(x_pointer == 4 && y_pointer == 8)
||(x_pointer == 155 && y_pointer == 8)
||(x_pointer == 156 && y_pointer == 8)
||(x_pointer == 157 && y_pointer == 8)
||(x_pointer == 2 && y_pointer == 9)
||(x_pointer == 3 && y_pointer == 9)
||(x_pointer == 4 && y_pointer == 9)
||(x_pointer == 155 && y_pointer == 9)
||(x_pointer == 156 && y_pointer == 9)
||(x_pointer == 157 && y_pointer == 9)
||(x_pointer == 2 && y_pointer == 10)
||(x_pointer == 3 && y_pointer == 10)
||(x_pointer == 4 && y_pointer == 10)
||(x_pointer == 155 && y_pointer == 10)
||(x_pointer == 156 && y_pointer == 10)
||(x_pointer == 157 && y_pointer == 10)
||(x_pointer == 2 && y_pointer == 11)
||(x_pointer == 3 && y_pointer == 11)
||(x_pointer == 4 && y_pointer == 11)
||(x_pointer == 155 && y_pointer == 11)
||(x_pointer == 156 && y_pointer == 11)
||(x_pointer == 157 && y_pointer == 11)
||(x_pointer == 2 && y_pointer == 12)
||(x_pointer == 3 && y_pointer == 12)
||(x_pointer == 4 && y_pointer == 12)
||(x_pointer == 155 && y_pointer == 12)
||(x_pointer == 156 && y_pointer == 12)
||(x_pointer == 157 && y_pointer == 12)
||(x_pointer == 2 && y_pointer == 13)
||(x_pointer == 3 && y_pointer == 13)
||(x_pointer == 4 && y_pointer == 13)
||(x_pointer == 155 && y_pointer == 13)
||(x_pointer == 156 && y_pointer == 13)
||(x_pointer == 157 && y_pointer == 13)
||(x_pointer == 2 && y_pointer == 14)
||(x_pointer == 3 && y_pointer == 14)
||(x_pointer == 4 && y_pointer == 14)
||(x_pointer == 14 && y_pointer == 14)
||(x_pointer == 15 && y_pointer == 14)
||(x_pointer == 16 && y_pointer == 14)
||(x_pointer == 17 && y_pointer == 14)
||(x_pointer == 18 && y_pointer == 14)
||(x_pointer == 19 && y_pointer == 14)
||(x_pointer == 20 && y_pointer == 14)
||(x_pointer == 21 && y_pointer == 14)
||(x_pointer == 22 && y_pointer == 14)
||(x_pointer == 32 && y_pointer == 14)
||(x_pointer == 33 && y_pointer == 14)
||(x_pointer == 34 && y_pointer == 14)
||(x_pointer == 35 && y_pointer == 14)
||(x_pointer == 36 && y_pointer == 14)
||(x_pointer == 37 && y_pointer == 14)
||(x_pointer == 38 && y_pointer == 14)
||(x_pointer == 39 && y_pointer == 14)
||(x_pointer == 40 && y_pointer == 14)
||(x_pointer == 50 && y_pointer == 14)
||(x_pointer == 51 && y_pointer == 14)
||(x_pointer == 52 && y_pointer == 14)
||(x_pointer == 53 && y_pointer == 14)
||(x_pointer == 54 && y_pointer == 14)
||(x_pointer == 55 && y_pointer == 14)
||(x_pointer == 56 && y_pointer == 14)
||(x_pointer == 57 && y_pointer == 14)
||(x_pointer == 58 && y_pointer == 14)
||(x_pointer == 68 && y_pointer == 14)
||(x_pointer == 69 && y_pointer == 14)
||(x_pointer == 70 && y_pointer == 14)
||(x_pointer == 71 && y_pointer == 14)
||(x_pointer == 72 && y_pointer == 14)
||(x_pointer == 73 && y_pointer == 14)
||(x_pointer == 74 && y_pointer == 14)
||(x_pointer == 75 && y_pointer == 14)
||(x_pointer == 76 && y_pointer == 14)
||(x_pointer == 86 && y_pointer == 14)
||(x_pointer == 87 && y_pointer == 14)
||(x_pointer == 88 && y_pointer == 14)
||(x_pointer == 89 && y_pointer == 14)
||(x_pointer == 90 && y_pointer == 14)
||(x_pointer == 91 && y_pointer == 14)
||(x_pointer == 92 && y_pointer == 14)
||(x_pointer == 93 && y_pointer == 14)
||(x_pointer == 94 && y_pointer == 14)
||(x_pointer == 104 && y_pointer == 14)
||(x_pointer == 105 && y_pointer == 14)
||(x_pointer == 106 && y_pointer == 14)
||(x_pointer == 107 && y_pointer == 14)
||(x_pointer == 108 && y_pointer == 14)
||(x_pointer == 109 && y_pointer == 14)
||(x_pointer == 110 && y_pointer == 14)
||(x_pointer == 111 && y_pointer == 14)
||(x_pointer == 112 && y_pointer == 14)
||(x_pointer == 122 && y_pointer == 14)
||(x_pointer == 123 && y_pointer == 14)
||(x_pointer == 124 && y_pointer == 14)
||(x_pointer == 125 && y_pointer == 14)
||(x_pointer == 126 && y_pointer == 14)
||(x_pointer == 127 && y_pointer == 14)
||(x_pointer == 128 && y_pointer == 14)
||(x_pointer == 129 && y_pointer == 14)
||(x_pointer == 130 && y_pointer == 14)
||(x_pointer == 140 && y_pointer == 14)
||(x_pointer == 141 && y_pointer == 14)
||(x_pointer == 142 && y_pointer == 14)
||(x_pointer == 143 && y_pointer == 14)
||(x_pointer == 144 && y_pointer == 14)
||(x_pointer == 145 && y_pointer == 14)
||(x_pointer == 146 && y_pointer == 14)
||(x_pointer == 147 && y_pointer == 14)
||(x_pointer == 148 && y_pointer == 14)
||(x_pointer == 155 && y_pointer == 14)
||(x_pointer == 156 && y_pointer == 14)
||(x_pointer == 157 && y_pointer == 14)
||(x_pointer == 2 && y_pointer == 15)
||(x_pointer == 3 && y_pointer == 15)
||(x_pointer == 4 && y_pointer == 15)
||(x_pointer == 14 && y_pointer == 15)
||(x_pointer == 15 && y_pointer == 15)
||(x_pointer == 16 && y_pointer == 15)
||(x_pointer == 17 && y_pointer == 15)
||(x_pointer == 18 && y_pointer == 15)
||(x_pointer == 19 && y_pointer == 15)
||(x_pointer == 20 && y_pointer == 15)
||(x_pointer == 21 && y_pointer == 15)
||(x_pointer == 22 && y_pointer == 15)
||(x_pointer == 32 && y_pointer == 15)
||(x_pointer == 33 && y_pointer == 15)
||(x_pointer == 34 && y_pointer == 15)
||(x_pointer == 35 && y_pointer == 15)
||(x_pointer == 36 && y_pointer == 15)
||(x_pointer == 37 && y_pointer == 15)
||(x_pointer == 38 && y_pointer == 15)
||(x_pointer == 39 && y_pointer == 15)
||(x_pointer == 40 && y_pointer == 15)
||(x_pointer == 50 && y_pointer == 15)
||(x_pointer == 51 && y_pointer == 15)
||(x_pointer == 52 && y_pointer == 15)
||(x_pointer == 53 && y_pointer == 15)
||(x_pointer == 54 && y_pointer == 15)
||(x_pointer == 55 && y_pointer == 15)
||(x_pointer == 56 && y_pointer == 15)
||(x_pointer == 57 && y_pointer == 15)
||(x_pointer == 58 && y_pointer == 15)
||(x_pointer == 68 && y_pointer == 15)
||(x_pointer == 69 && y_pointer == 15)
||(x_pointer == 70 && y_pointer == 15)
||(x_pointer == 71 && y_pointer == 15)
||(x_pointer == 72 && y_pointer == 15)
||(x_pointer == 73 && y_pointer == 15)
||(x_pointer == 74 && y_pointer == 15)
||(x_pointer == 75 && y_pointer == 15)
||(x_pointer == 76 && y_pointer == 15)
||(x_pointer == 86 && y_pointer == 15)
||(x_pointer == 87 && y_pointer == 15)
||(x_pointer == 88 && y_pointer == 15)
||(x_pointer == 89 && y_pointer == 15)
||(x_pointer == 90 && y_pointer == 15)
||(x_pointer == 91 && y_pointer == 15)
||(x_pointer == 92 && y_pointer == 15)
||(x_pointer == 93 && y_pointer == 15)
||(x_pointer == 94 && y_pointer == 15)
||(x_pointer == 104 && y_pointer == 15)
||(x_pointer == 105 && y_pointer == 15)
||(x_pointer == 106 && y_pointer == 15)
||(x_pointer == 107 && y_pointer == 15)
||(x_pointer == 108 && y_pointer == 15)
||(x_pointer == 109 && y_pointer == 15)
||(x_pointer == 110 && y_pointer == 15)
||(x_pointer == 111 && y_pointer == 15)
||(x_pointer == 112 && y_pointer == 15)
||(x_pointer == 122 && y_pointer == 15)
||(x_pointer == 123 && y_pointer == 15)
||(x_pointer == 124 && y_pointer == 15)
||(x_pointer == 125 && y_pointer == 15)
||(x_pointer == 126 && y_pointer == 15)
||(x_pointer == 127 && y_pointer == 15)
||(x_pointer == 128 && y_pointer == 15)
||(x_pointer == 129 && y_pointer == 15)
||(x_pointer == 130 && y_pointer == 15)
||(x_pointer == 140 && y_pointer == 15)
||(x_pointer == 141 && y_pointer == 15)
||(x_pointer == 142 && y_pointer == 15)
||(x_pointer == 143 && y_pointer == 15)
||(x_pointer == 144 && y_pointer == 15)
||(x_pointer == 145 && y_pointer == 15)
||(x_pointer == 146 && y_pointer == 15)
||(x_pointer == 147 && y_pointer == 15)
||(x_pointer == 148 && y_pointer == 15)
||(x_pointer == 155 && y_pointer == 15)
||(x_pointer == 156 && y_pointer == 15)
||(x_pointer == 157 && y_pointer == 15)
||(x_pointer == 2 && y_pointer == 16)
||(x_pointer == 3 && y_pointer == 16)
||(x_pointer == 4 && y_pointer == 16)
||(x_pointer == 14 && y_pointer == 16)
||(x_pointer == 15 && y_pointer == 16)
||(x_pointer == 16 && y_pointer == 16)
||(x_pointer == 17 && y_pointer == 16)
||(x_pointer == 18 && y_pointer == 16)
||(x_pointer == 19 && y_pointer == 16)
||(x_pointer == 20 && y_pointer == 16)
||(x_pointer == 21 && y_pointer == 16)
||(x_pointer == 22 && y_pointer == 16)
||(x_pointer == 32 && y_pointer == 16)
||(x_pointer == 33 && y_pointer == 16)
||(x_pointer == 34 && y_pointer == 16)
||(x_pointer == 35 && y_pointer == 16)
||(x_pointer == 36 && y_pointer == 16)
||(x_pointer == 37 && y_pointer == 16)
||(x_pointer == 38 && y_pointer == 16)
||(x_pointer == 39 && y_pointer == 16)
||(x_pointer == 40 && y_pointer == 16)
||(x_pointer == 50 && y_pointer == 16)
||(x_pointer == 51 && y_pointer == 16)
||(x_pointer == 52 && y_pointer == 16)
||(x_pointer == 53 && y_pointer == 16)
||(x_pointer == 54 && y_pointer == 16)
||(x_pointer == 55 && y_pointer == 16)
||(x_pointer == 56 && y_pointer == 16)
||(x_pointer == 57 && y_pointer == 16)
||(x_pointer == 58 && y_pointer == 16)
||(x_pointer == 68 && y_pointer == 16)
||(x_pointer == 69 && y_pointer == 16)
||(x_pointer == 70 && y_pointer == 16)
||(x_pointer == 71 && y_pointer == 16)
||(x_pointer == 72 && y_pointer == 16)
||(x_pointer == 73 && y_pointer == 16)
||(x_pointer == 74 && y_pointer == 16)
||(x_pointer == 75 && y_pointer == 16)
||(x_pointer == 76 && y_pointer == 16)
||(x_pointer == 86 && y_pointer == 16)
||(x_pointer == 87 && y_pointer == 16)
||(x_pointer == 88 && y_pointer == 16)
||(x_pointer == 89 && y_pointer == 16)
||(x_pointer == 90 && y_pointer == 16)
||(x_pointer == 91 && y_pointer == 16)
||(x_pointer == 92 && y_pointer == 16)
||(x_pointer == 93 && y_pointer == 16)
||(x_pointer == 94 && y_pointer == 16)
||(x_pointer == 104 && y_pointer == 16)
||(x_pointer == 105 && y_pointer == 16)
||(x_pointer == 106 && y_pointer == 16)
||(x_pointer == 107 && y_pointer == 16)
||(x_pointer == 108 && y_pointer == 16)
||(x_pointer == 109 && y_pointer == 16)
||(x_pointer == 110 && y_pointer == 16)
||(x_pointer == 111 && y_pointer == 16)
||(x_pointer == 112 && y_pointer == 16)
||(x_pointer == 122 && y_pointer == 16)
||(x_pointer == 123 && y_pointer == 16)
||(x_pointer == 124 && y_pointer == 16)
||(x_pointer == 125 && y_pointer == 16)
||(x_pointer == 126 && y_pointer == 16)
||(x_pointer == 127 && y_pointer == 16)
||(x_pointer == 128 && y_pointer == 16)
||(x_pointer == 129 && y_pointer == 16)
||(x_pointer == 130 && y_pointer == 16)
||(x_pointer == 140 && y_pointer == 16)
||(x_pointer == 141 && y_pointer == 16)
||(x_pointer == 142 && y_pointer == 16)
||(x_pointer == 143 && y_pointer == 16)
||(x_pointer == 144 && y_pointer == 16)
||(x_pointer == 145 && y_pointer == 16)
||(x_pointer == 146 && y_pointer == 16)
||(x_pointer == 147 && y_pointer == 16)
||(x_pointer == 148 && y_pointer == 16)
||(x_pointer == 155 && y_pointer == 16)
||(x_pointer == 156 && y_pointer == 16)
||(x_pointer == 157 && y_pointer == 16)
||(x_pointer == 2 && y_pointer == 17)
||(x_pointer == 3 && y_pointer == 17)
||(x_pointer == 4 && y_pointer == 17)
||(x_pointer == 14 && y_pointer == 17)
||(x_pointer == 15 && y_pointer == 17)
||(x_pointer == 16 && y_pointer == 17)
||(x_pointer == 17 && y_pointer == 17)
||(x_pointer == 18 && y_pointer == 17)
||(x_pointer == 19 && y_pointer == 17)
||(x_pointer == 20 && y_pointer == 17)
||(x_pointer == 21 && y_pointer == 17)
||(x_pointer == 22 && y_pointer == 17)
||(x_pointer == 32 && y_pointer == 17)
||(x_pointer == 33 && y_pointer == 17)
||(x_pointer == 34 && y_pointer == 17)
||(x_pointer == 35 && y_pointer == 17)
||(x_pointer == 36 && y_pointer == 17)
||(x_pointer == 37 && y_pointer == 17)
||(x_pointer == 38 && y_pointer == 17)
||(x_pointer == 39 && y_pointer == 17)
||(x_pointer == 40 && y_pointer == 17)
||(x_pointer == 50 && y_pointer == 17)
||(x_pointer == 51 && y_pointer == 17)
||(x_pointer == 52 && y_pointer == 17)
||(x_pointer == 53 && y_pointer == 17)
||(x_pointer == 54 && y_pointer == 17)
||(x_pointer == 55 && y_pointer == 17)
||(x_pointer == 56 && y_pointer == 17)
||(x_pointer == 57 && y_pointer == 17)
||(x_pointer == 58 && y_pointer == 17)
||(x_pointer == 68 && y_pointer == 17)
||(x_pointer == 69 && y_pointer == 17)
||(x_pointer == 70 && y_pointer == 17)
||(x_pointer == 71 && y_pointer == 17)
||(x_pointer == 72 && y_pointer == 17)
||(x_pointer == 73 && y_pointer == 17)
||(x_pointer == 74 && y_pointer == 17)
||(x_pointer == 75 && y_pointer == 17)
||(x_pointer == 76 && y_pointer == 17)
||(x_pointer == 86 && y_pointer == 17)
||(x_pointer == 87 && y_pointer == 17)
||(x_pointer == 88 && y_pointer == 17)
||(x_pointer == 89 && y_pointer == 17)
||(x_pointer == 90 && y_pointer == 17)
||(x_pointer == 91 && y_pointer == 17)
||(x_pointer == 92 && y_pointer == 17)
||(x_pointer == 93 && y_pointer == 17)
||(x_pointer == 94 && y_pointer == 17)
||(x_pointer == 104 && y_pointer == 17)
||(x_pointer == 105 && y_pointer == 17)
||(x_pointer == 106 && y_pointer == 17)
||(x_pointer == 107 && y_pointer == 17)
||(x_pointer == 108 && y_pointer == 17)
||(x_pointer == 109 && y_pointer == 17)
||(x_pointer == 110 && y_pointer == 17)
||(x_pointer == 111 && y_pointer == 17)
||(x_pointer == 112 && y_pointer == 17)
||(x_pointer == 122 && y_pointer == 17)
||(x_pointer == 123 && y_pointer == 17)
||(x_pointer == 124 && y_pointer == 17)
||(x_pointer == 125 && y_pointer == 17)
||(x_pointer == 126 && y_pointer == 17)
||(x_pointer == 127 && y_pointer == 17)
||(x_pointer == 128 && y_pointer == 17)
||(x_pointer == 129 && y_pointer == 17)
||(x_pointer == 130 && y_pointer == 17)
||(x_pointer == 140 && y_pointer == 17)
||(x_pointer == 141 && y_pointer == 17)
||(x_pointer == 142 && y_pointer == 17)
||(x_pointer == 143 && y_pointer == 17)
||(x_pointer == 144 && y_pointer == 17)
||(x_pointer == 145 && y_pointer == 17)
||(x_pointer == 146 && y_pointer == 17)
||(x_pointer == 147 && y_pointer == 17)
||(x_pointer == 148 && y_pointer == 17)
||(x_pointer == 155 && y_pointer == 17)
||(x_pointer == 156 && y_pointer == 17)
||(x_pointer == 157 && y_pointer == 17)
||(x_pointer == 2 && y_pointer == 18)
||(x_pointer == 3 && y_pointer == 18)
||(x_pointer == 4 && y_pointer == 18)
||(x_pointer == 14 && y_pointer == 18)
||(x_pointer == 15 && y_pointer == 18)
||(x_pointer == 16 && y_pointer == 18)
||(x_pointer == 17 && y_pointer == 18)
||(x_pointer == 18 && y_pointer == 18)
||(x_pointer == 19 && y_pointer == 18)
||(x_pointer == 20 && y_pointer == 18)
||(x_pointer == 21 && y_pointer == 18)
||(x_pointer == 22 && y_pointer == 18)
||(x_pointer == 32 && y_pointer == 18)
||(x_pointer == 33 && y_pointer == 18)
||(x_pointer == 34 && y_pointer == 18)
||(x_pointer == 35 && y_pointer == 18)
||(x_pointer == 36 && y_pointer == 18)
||(x_pointer == 37 && y_pointer == 18)
||(x_pointer == 38 && y_pointer == 18)
||(x_pointer == 39 && y_pointer == 18)
||(x_pointer == 40 && y_pointer == 18)
||(x_pointer == 50 && y_pointer == 18)
||(x_pointer == 51 && y_pointer == 18)
||(x_pointer == 52 && y_pointer == 18)
||(x_pointer == 53 && y_pointer == 18)
||(x_pointer == 54 && y_pointer == 18)
||(x_pointer == 55 && y_pointer == 18)
||(x_pointer == 56 && y_pointer == 18)
||(x_pointer == 57 && y_pointer == 18)
||(x_pointer == 58 && y_pointer == 18)
||(x_pointer == 68 && y_pointer == 18)
||(x_pointer == 69 && y_pointer == 18)
||(x_pointer == 70 && y_pointer == 18)
||(x_pointer == 71 && y_pointer == 18)
||(x_pointer == 72 && y_pointer == 18)
||(x_pointer == 73 && y_pointer == 18)
||(x_pointer == 74 && y_pointer == 18)
||(x_pointer == 75 && y_pointer == 18)
||(x_pointer == 76 && y_pointer == 18)
||(x_pointer == 86 && y_pointer == 18)
||(x_pointer == 87 && y_pointer == 18)
||(x_pointer == 88 && y_pointer == 18)
||(x_pointer == 89 && y_pointer == 18)
||(x_pointer == 90 && y_pointer == 18)
||(x_pointer == 91 && y_pointer == 18)
||(x_pointer == 92 && y_pointer == 18)
||(x_pointer == 93 && y_pointer == 18)
||(x_pointer == 94 && y_pointer == 18)
||(x_pointer == 104 && y_pointer == 18)
||(x_pointer == 105 && y_pointer == 18)
||(x_pointer == 106 && y_pointer == 18)
||(x_pointer == 107 && y_pointer == 18)
||(x_pointer == 108 && y_pointer == 18)
||(x_pointer == 109 && y_pointer == 18)
||(x_pointer == 110 && y_pointer == 18)
||(x_pointer == 111 && y_pointer == 18)
||(x_pointer == 112 && y_pointer == 18)
||(x_pointer == 122 && y_pointer == 18)
||(x_pointer == 123 && y_pointer == 18)
||(x_pointer == 124 && y_pointer == 18)
||(x_pointer == 125 && y_pointer == 18)
||(x_pointer == 126 && y_pointer == 18)
||(x_pointer == 127 && y_pointer == 18)
||(x_pointer == 128 && y_pointer == 18)
||(x_pointer == 129 && y_pointer == 18)
||(x_pointer == 130 && y_pointer == 18)
||(x_pointer == 140 && y_pointer == 18)
||(x_pointer == 141 && y_pointer == 18)
||(x_pointer == 142 && y_pointer == 18)
||(x_pointer == 143 && y_pointer == 18)
||(x_pointer == 144 && y_pointer == 18)
||(x_pointer == 145 && y_pointer == 18)
||(x_pointer == 146 && y_pointer == 18)
||(x_pointer == 147 && y_pointer == 18)
||(x_pointer == 148 && y_pointer == 18)
||(x_pointer == 155 && y_pointer == 18)
||(x_pointer == 156 && y_pointer == 18)
||(x_pointer == 157 && y_pointer == 18)
||(x_pointer == 2 && y_pointer == 19)
||(x_pointer == 3 && y_pointer == 19)
||(x_pointer == 4 && y_pointer == 19)
||(x_pointer == 14 && y_pointer == 19)
||(x_pointer == 15 && y_pointer == 19)
||(x_pointer == 16 && y_pointer == 19)
||(x_pointer == 17 && y_pointer == 19)
||(x_pointer == 18 && y_pointer == 19)
||(x_pointer == 19 && y_pointer == 19)
||(x_pointer == 20 && y_pointer == 19)
||(x_pointer == 21 && y_pointer == 19)
||(x_pointer == 22 && y_pointer == 19)
||(x_pointer == 32 && y_pointer == 19)
||(x_pointer == 33 && y_pointer == 19)
||(x_pointer == 34 && y_pointer == 19)
||(x_pointer == 35 && y_pointer == 19)
||(x_pointer == 36 && y_pointer == 19)
||(x_pointer == 37 && y_pointer == 19)
||(x_pointer == 38 && y_pointer == 19)
||(x_pointer == 39 && y_pointer == 19)
||(x_pointer == 40 && y_pointer == 19)
||(x_pointer == 50 && y_pointer == 19)
||(x_pointer == 51 && y_pointer == 19)
||(x_pointer == 52 && y_pointer == 19)
||(x_pointer == 53 && y_pointer == 19)
||(x_pointer == 54 && y_pointer == 19)
||(x_pointer == 55 && y_pointer == 19)
||(x_pointer == 56 && y_pointer == 19)
||(x_pointer == 57 && y_pointer == 19)
||(x_pointer == 58 && y_pointer == 19)
||(x_pointer == 68 && y_pointer == 19)
||(x_pointer == 69 && y_pointer == 19)
||(x_pointer == 70 && y_pointer == 19)
||(x_pointer == 71 && y_pointer == 19)
||(x_pointer == 72 && y_pointer == 19)
||(x_pointer == 73 && y_pointer == 19)
||(x_pointer == 74 && y_pointer == 19)
||(x_pointer == 75 && y_pointer == 19)
||(x_pointer == 76 && y_pointer == 19)
||(x_pointer == 86 && y_pointer == 19)
||(x_pointer == 87 && y_pointer == 19)
||(x_pointer == 88 && y_pointer == 19)
||(x_pointer == 89 && y_pointer == 19)
||(x_pointer == 90 && y_pointer == 19)
||(x_pointer == 91 && y_pointer == 19)
||(x_pointer == 92 && y_pointer == 19)
||(x_pointer == 93 && y_pointer == 19)
||(x_pointer == 94 && y_pointer == 19)
||(x_pointer == 104 && y_pointer == 19)
||(x_pointer == 105 && y_pointer == 19)
||(x_pointer == 106 && y_pointer == 19)
||(x_pointer == 107 && y_pointer == 19)
||(x_pointer == 108 && y_pointer == 19)
||(x_pointer == 109 && y_pointer == 19)
||(x_pointer == 110 && y_pointer == 19)
||(x_pointer == 111 && y_pointer == 19)
||(x_pointer == 112 && y_pointer == 19)
||(x_pointer == 122 && y_pointer == 19)
||(x_pointer == 123 && y_pointer == 19)
||(x_pointer == 124 && y_pointer == 19)
||(x_pointer == 125 && y_pointer == 19)
||(x_pointer == 126 && y_pointer == 19)
||(x_pointer == 127 && y_pointer == 19)
||(x_pointer == 128 && y_pointer == 19)
||(x_pointer == 129 && y_pointer == 19)
||(x_pointer == 130 && y_pointer == 19)
||(x_pointer == 140 && y_pointer == 19)
||(x_pointer == 141 && y_pointer == 19)
||(x_pointer == 142 && y_pointer == 19)
||(x_pointer == 143 && y_pointer == 19)
||(x_pointer == 144 && y_pointer == 19)
||(x_pointer == 145 && y_pointer == 19)
||(x_pointer == 146 && y_pointer == 19)
||(x_pointer == 147 && y_pointer == 19)
||(x_pointer == 148 && y_pointer == 19)
||(x_pointer == 155 && y_pointer == 19)
||(x_pointer == 156 && y_pointer == 19)
||(x_pointer == 157 && y_pointer == 19)
||(x_pointer == 2 && y_pointer == 20)
||(x_pointer == 3 && y_pointer == 20)
||(x_pointer == 4 && y_pointer == 20)
||(x_pointer == 14 && y_pointer == 20)
||(x_pointer == 15 && y_pointer == 20)
||(x_pointer == 16 && y_pointer == 20)
||(x_pointer == 17 && y_pointer == 20)
||(x_pointer == 18 && y_pointer == 20)
||(x_pointer == 19 && y_pointer == 20)
||(x_pointer == 20 && y_pointer == 20)
||(x_pointer == 21 && y_pointer == 20)
||(x_pointer == 22 && y_pointer == 20)
||(x_pointer == 32 && y_pointer == 20)
||(x_pointer == 33 && y_pointer == 20)
||(x_pointer == 34 && y_pointer == 20)
||(x_pointer == 35 && y_pointer == 20)
||(x_pointer == 36 && y_pointer == 20)
||(x_pointer == 37 && y_pointer == 20)
||(x_pointer == 38 && y_pointer == 20)
||(x_pointer == 39 && y_pointer == 20)
||(x_pointer == 40 && y_pointer == 20)
||(x_pointer == 50 && y_pointer == 20)
||(x_pointer == 51 && y_pointer == 20)
||(x_pointer == 52 && y_pointer == 20)
||(x_pointer == 53 && y_pointer == 20)
||(x_pointer == 54 && y_pointer == 20)
||(x_pointer == 55 && y_pointer == 20)
||(x_pointer == 56 && y_pointer == 20)
||(x_pointer == 57 && y_pointer == 20)
||(x_pointer == 58 && y_pointer == 20)
||(x_pointer == 68 && y_pointer == 20)
||(x_pointer == 69 && y_pointer == 20)
||(x_pointer == 70 && y_pointer == 20)
||(x_pointer == 71 && y_pointer == 20)
||(x_pointer == 72 && y_pointer == 20)
||(x_pointer == 73 && y_pointer == 20)
||(x_pointer == 74 && y_pointer == 20)
||(x_pointer == 75 && y_pointer == 20)
||(x_pointer == 76 && y_pointer == 20)
||(x_pointer == 86 && y_pointer == 20)
||(x_pointer == 87 && y_pointer == 20)
||(x_pointer == 88 && y_pointer == 20)
||(x_pointer == 89 && y_pointer == 20)
||(x_pointer == 90 && y_pointer == 20)
||(x_pointer == 91 && y_pointer == 20)
||(x_pointer == 92 && y_pointer == 20)
||(x_pointer == 93 && y_pointer == 20)
||(x_pointer == 94 && y_pointer == 20)
||(x_pointer == 104 && y_pointer == 20)
||(x_pointer == 105 && y_pointer == 20)
||(x_pointer == 106 && y_pointer == 20)
||(x_pointer == 107 && y_pointer == 20)
||(x_pointer == 108 && y_pointer == 20)
||(x_pointer == 109 && y_pointer == 20)
||(x_pointer == 110 && y_pointer == 20)
||(x_pointer == 111 && y_pointer == 20)
||(x_pointer == 112 && y_pointer == 20)
||(x_pointer == 122 && y_pointer == 20)
||(x_pointer == 123 && y_pointer == 20)
||(x_pointer == 124 && y_pointer == 20)
||(x_pointer == 125 && y_pointer == 20)
||(x_pointer == 126 && y_pointer == 20)
||(x_pointer == 127 && y_pointer == 20)
||(x_pointer == 128 && y_pointer == 20)
||(x_pointer == 129 && y_pointer == 20)
||(x_pointer == 130 && y_pointer == 20)
||(x_pointer == 140 && y_pointer == 20)
||(x_pointer == 141 && y_pointer == 20)
||(x_pointer == 142 && y_pointer == 20)
||(x_pointer == 143 && y_pointer == 20)
||(x_pointer == 144 && y_pointer == 20)
||(x_pointer == 145 && y_pointer == 20)
||(x_pointer == 146 && y_pointer == 20)
||(x_pointer == 147 && y_pointer == 20)
||(x_pointer == 148 && y_pointer == 20)
||(x_pointer == 155 && y_pointer == 20)
||(x_pointer == 156 && y_pointer == 20)
||(x_pointer == 157 && y_pointer == 20)
||(x_pointer == 2 && y_pointer == 21)
||(x_pointer == 3 && y_pointer == 21)
||(x_pointer == 4 && y_pointer == 21)
||(x_pointer == 14 && y_pointer == 21)
||(x_pointer == 15 && y_pointer == 21)
||(x_pointer == 16 && y_pointer == 21)
||(x_pointer == 17 && y_pointer == 21)
||(x_pointer == 18 && y_pointer == 21)
||(x_pointer == 19 && y_pointer == 21)
||(x_pointer == 20 && y_pointer == 21)
||(x_pointer == 21 && y_pointer == 21)
||(x_pointer == 22 && y_pointer == 21)
||(x_pointer == 32 && y_pointer == 21)
||(x_pointer == 33 && y_pointer == 21)
||(x_pointer == 34 && y_pointer == 21)
||(x_pointer == 35 && y_pointer == 21)
||(x_pointer == 36 && y_pointer == 21)
||(x_pointer == 37 && y_pointer == 21)
||(x_pointer == 38 && y_pointer == 21)
||(x_pointer == 39 && y_pointer == 21)
||(x_pointer == 40 && y_pointer == 21)
||(x_pointer == 50 && y_pointer == 21)
||(x_pointer == 51 && y_pointer == 21)
||(x_pointer == 52 && y_pointer == 21)
||(x_pointer == 53 && y_pointer == 21)
||(x_pointer == 54 && y_pointer == 21)
||(x_pointer == 55 && y_pointer == 21)
||(x_pointer == 56 && y_pointer == 21)
||(x_pointer == 57 && y_pointer == 21)
||(x_pointer == 58 && y_pointer == 21)
||(x_pointer == 68 && y_pointer == 21)
||(x_pointer == 69 && y_pointer == 21)
||(x_pointer == 70 && y_pointer == 21)
||(x_pointer == 71 && y_pointer == 21)
||(x_pointer == 72 && y_pointer == 21)
||(x_pointer == 73 && y_pointer == 21)
||(x_pointer == 74 && y_pointer == 21)
||(x_pointer == 75 && y_pointer == 21)
||(x_pointer == 76 && y_pointer == 21)
||(x_pointer == 86 && y_pointer == 21)
||(x_pointer == 87 && y_pointer == 21)
||(x_pointer == 88 && y_pointer == 21)
||(x_pointer == 89 && y_pointer == 21)
||(x_pointer == 90 && y_pointer == 21)
||(x_pointer == 91 && y_pointer == 21)
||(x_pointer == 92 && y_pointer == 21)
||(x_pointer == 93 && y_pointer == 21)
||(x_pointer == 94 && y_pointer == 21)
||(x_pointer == 104 && y_pointer == 21)
||(x_pointer == 105 && y_pointer == 21)
||(x_pointer == 106 && y_pointer == 21)
||(x_pointer == 107 && y_pointer == 21)
||(x_pointer == 108 && y_pointer == 21)
||(x_pointer == 109 && y_pointer == 21)
||(x_pointer == 110 && y_pointer == 21)
||(x_pointer == 111 && y_pointer == 21)
||(x_pointer == 112 && y_pointer == 21)
||(x_pointer == 122 && y_pointer == 21)
||(x_pointer == 123 && y_pointer == 21)
||(x_pointer == 124 && y_pointer == 21)
||(x_pointer == 125 && y_pointer == 21)
||(x_pointer == 126 && y_pointer == 21)
||(x_pointer == 127 && y_pointer == 21)
||(x_pointer == 128 && y_pointer == 21)
||(x_pointer == 129 && y_pointer == 21)
||(x_pointer == 130 && y_pointer == 21)
||(x_pointer == 140 && y_pointer == 21)
||(x_pointer == 141 && y_pointer == 21)
||(x_pointer == 142 && y_pointer == 21)
||(x_pointer == 143 && y_pointer == 21)
||(x_pointer == 144 && y_pointer == 21)
||(x_pointer == 145 && y_pointer == 21)
||(x_pointer == 146 && y_pointer == 21)
||(x_pointer == 147 && y_pointer == 21)
||(x_pointer == 148 && y_pointer == 21)
||(x_pointer == 155 && y_pointer == 21)
||(x_pointer == 156 && y_pointer == 21)
||(x_pointer == 157 && y_pointer == 21)
||(x_pointer == 2 && y_pointer == 22)
||(x_pointer == 3 && y_pointer == 22)
||(x_pointer == 4 && y_pointer == 22)
||(x_pointer == 14 && y_pointer == 22)
||(x_pointer == 15 && y_pointer == 22)
||(x_pointer == 16 && y_pointer == 22)
||(x_pointer == 17 && y_pointer == 22)
||(x_pointer == 18 && y_pointer == 22)
||(x_pointer == 19 && y_pointer == 22)
||(x_pointer == 20 && y_pointer == 22)
||(x_pointer == 21 && y_pointer == 22)
||(x_pointer == 22 && y_pointer == 22)
||(x_pointer == 32 && y_pointer == 22)
||(x_pointer == 33 && y_pointer == 22)
||(x_pointer == 34 && y_pointer == 22)
||(x_pointer == 35 && y_pointer == 22)
||(x_pointer == 36 && y_pointer == 22)
||(x_pointer == 37 && y_pointer == 22)
||(x_pointer == 38 && y_pointer == 22)
||(x_pointer == 39 && y_pointer == 22)
||(x_pointer == 40 && y_pointer == 22)
||(x_pointer == 50 && y_pointer == 22)
||(x_pointer == 51 && y_pointer == 22)
||(x_pointer == 52 && y_pointer == 22)
||(x_pointer == 53 && y_pointer == 22)
||(x_pointer == 54 && y_pointer == 22)
||(x_pointer == 55 && y_pointer == 22)
||(x_pointer == 56 && y_pointer == 22)
||(x_pointer == 57 && y_pointer == 22)
||(x_pointer == 58 && y_pointer == 22)
||(x_pointer == 68 && y_pointer == 22)
||(x_pointer == 69 && y_pointer == 22)
||(x_pointer == 70 && y_pointer == 22)
||(x_pointer == 71 && y_pointer == 22)
||(x_pointer == 72 && y_pointer == 22)
||(x_pointer == 73 && y_pointer == 22)
||(x_pointer == 74 && y_pointer == 22)
||(x_pointer == 75 && y_pointer == 22)
||(x_pointer == 76 && y_pointer == 22)
||(x_pointer == 86 && y_pointer == 22)
||(x_pointer == 87 && y_pointer == 22)
||(x_pointer == 88 && y_pointer == 22)
||(x_pointer == 89 && y_pointer == 22)
||(x_pointer == 90 && y_pointer == 22)
||(x_pointer == 91 && y_pointer == 22)
||(x_pointer == 92 && y_pointer == 22)
||(x_pointer == 93 && y_pointer == 22)
||(x_pointer == 94 && y_pointer == 22)
||(x_pointer == 104 && y_pointer == 22)
||(x_pointer == 105 && y_pointer == 22)
||(x_pointer == 106 && y_pointer == 22)
||(x_pointer == 107 && y_pointer == 22)
||(x_pointer == 108 && y_pointer == 22)
||(x_pointer == 109 && y_pointer == 22)
||(x_pointer == 110 && y_pointer == 22)
||(x_pointer == 111 && y_pointer == 22)
||(x_pointer == 112 && y_pointer == 22)
||(x_pointer == 122 && y_pointer == 22)
||(x_pointer == 123 && y_pointer == 22)
||(x_pointer == 124 && y_pointer == 22)
||(x_pointer == 125 && y_pointer == 22)
||(x_pointer == 126 && y_pointer == 22)
||(x_pointer == 127 && y_pointer == 22)
||(x_pointer == 128 && y_pointer == 22)
||(x_pointer == 129 && y_pointer == 22)
||(x_pointer == 130 && y_pointer == 22)
||(x_pointer == 140 && y_pointer == 22)
||(x_pointer == 141 && y_pointer == 22)
||(x_pointer == 142 && y_pointer == 22)
||(x_pointer == 143 && y_pointer == 22)
||(x_pointer == 144 && y_pointer == 22)
||(x_pointer == 145 && y_pointer == 22)
||(x_pointer == 146 && y_pointer == 22)
||(x_pointer == 147 && y_pointer == 22)
||(x_pointer == 148 && y_pointer == 22)
||(x_pointer == 155 && y_pointer == 22)
||(x_pointer == 156 && y_pointer == 22)
||(x_pointer == 157 && y_pointer == 22)
||(x_pointer == 2 && y_pointer == 23)
||(x_pointer == 3 && y_pointer == 23)
||(x_pointer == 4 && y_pointer == 23)
||(x_pointer == 155 && y_pointer == 23)
||(x_pointer == 156 && y_pointer == 23)
||(x_pointer == 157 && y_pointer == 23)
||(x_pointer == 2 && y_pointer == 24)
||(x_pointer == 3 && y_pointer == 24)
||(x_pointer == 4 && y_pointer == 24)
||(x_pointer == 155 && y_pointer == 24)
||(x_pointer == 156 && y_pointer == 24)
||(x_pointer == 157 && y_pointer == 24)
||(x_pointer == 2 && y_pointer == 25)
||(x_pointer == 3 && y_pointer == 25)
||(x_pointer == 4 && y_pointer == 25)
||(x_pointer == 155 && y_pointer == 25)
||(x_pointer == 156 && y_pointer == 25)
||(x_pointer == 157 && y_pointer == 25)
||(x_pointer == 2 && y_pointer == 26)
||(x_pointer == 3 && y_pointer == 26)
||(x_pointer == 4 && y_pointer == 26)
||(x_pointer == 155 && y_pointer == 26)
||(x_pointer == 156 && y_pointer == 26)
||(x_pointer == 157 && y_pointer == 26)
||(x_pointer == 2 && y_pointer == 27)
||(x_pointer == 3 && y_pointer == 27)
||(x_pointer == 4 && y_pointer == 27)
||(x_pointer == 155 && y_pointer == 27)
||(x_pointer == 156 && y_pointer == 27)
||(x_pointer == 157 && y_pointer == 27)
||(x_pointer == 2 && y_pointer == 28)
||(x_pointer == 3 && y_pointer == 28)
||(x_pointer == 4 && y_pointer == 28)
||(x_pointer == 155 && y_pointer == 28)
||(x_pointer == 156 && y_pointer == 28)
||(x_pointer == 157 && y_pointer == 28)
||(x_pointer == 2 && y_pointer == 29)
||(x_pointer == 3 && y_pointer == 29)
||(x_pointer == 4 && y_pointer == 29)
||(x_pointer == 155 && y_pointer == 29)
||(x_pointer == 156 && y_pointer == 29)
||(x_pointer == 157 && y_pointer == 29)
||(x_pointer == 2 && y_pointer == 30)
||(x_pointer == 3 && y_pointer == 30)
||(x_pointer == 4 && y_pointer == 30)
||(x_pointer == 155 && y_pointer == 30)
||(x_pointer == 156 && y_pointer == 30)
||(x_pointer == 157 && y_pointer == 30)
||(x_pointer == 2 && y_pointer == 31)
||(x_pointer == 3 && y_pointer == 31)
||(x_pointer == 4 && y_pointer == 31)
||(x_pointer == 155 && y_pointer == 31)
||(x_pointer == 156 && y_pointer == 31)
||(x_pointer == 157 && y_pointer == 31)
||(x_pointer == 2 && y_pointer == 32)
||(x_pointer == 3 && y_pointer == 32)
||(x_pointer == 4 && y_pointer == 32)
||(x_pointer == 14 && y_pointer == 32)
||(x_pointer == 15 && y_pointer == 32)
||(x_pointer == 16 && y_pointer == 32)
||(x_pointer == 17 && y_pointer == 32)
||(x_pointer == 18 && y_pointer == 32)
||(x_pointer == 19 && y_pointer == 32)
||(x_pointer == 20 && y_pointer == 32)
||(x_pointer == 21 && y_pointer == 32)
||(x_pointer == 22 && y_pointer == 32)
||(x_pointer == 32 && y_pointer == 32)
||(x_pointer == 33 && y_pointer == 32)
||(x_pointer == 34 && y_pointer == 32)
||(x_pointer == 35 && y_pointer == 32)
||(x_pointer == 36 && y_pointer == 32)
||(x_pointer == 37 && y_pointer == 32)
||(x_pointer == 38 && y_pointer == 32)
||(x_pointer == 39 && y_pointer == 32)
||(x_pointer == 40 && y_pointer == 32)
||(x_pointer == 50 && y_pointer == 32)
||(x_pointer == 51 && y_pointer == 32)
||(x_pointer == 52 && y_pointer == 32)
||(x_pointer == 53 && y_pointer == 32)
||(x_pointer == 54 && y_pointer == 32)
||(x_pointer == 55 && y_pointer == 32)
||(x_pointer == 56 && y_pointer == 32)
||(x_pointer == 57 && y_pointer == 32)
||(x_pointer == 58 && y_pointer == 32)
||(x_pointer == 68 && y_pointer == 32)
||(x_pointer == 69 && y_pointer == 32)
||(x_pointer == 70 && y_pointer == 32)
||(x_pointer == 71 && y_pointer == 32)
||(x_pointer == 72 && y_pointer == 32)
||(x_pointer == 73 && y_pointer == 32)
||(x_pointer == 74 && y_pointer == 32)
||(x_pointer == 75 && y_pointer == 32)
||(x_pointer == 76 && y_pointer == 32)
||(x_pointer == 86 && y_pointer == 32)
||(x_pointer == 87 && y_pointer == 32)
||(x_pointer == 88 && y_pointer == 32)
||(x_pointer == 89 && y_pointer == 32)
||(x_pointer == 90 && y_pointer == 32)
||(x_pointer == 91 && y_pointer == 32)
||(x_pointer == 92 && y_pointer == 32)
||(x_pointer == 93 && y_pointer == 32)
||(x_pointer == 94 && y_pointer == 32)
||(x_pointer == 104 && y_pointer == 32)
||(x_pointer == 105 && y_pointer == 32)
||(x_pointer == 106 && y_pointer == 32)
||(x_pointer == 107 && y_pointer == 32)
||(x_pointer == 108 && y_pointer == 32)
||(x_pointer == 109 && y_pointer == 32)
||(x_pointer == 110 && y_pointer == 32)
||(x_pointer == 111 && y_pointer == 32)
||(x_pointer == 112 && y_pointer == 32)
||(x_pointer == 122 && y_pointer == 32)
||(x_pointer == 123 && y_pointer == 32)
||(x_pointer == 124 && y_pointer == 32)
||(x_pointer == 125 && y_pointer == 32)
||(x_pointer == 126 && y_pointer == 32)
||(x_pointer == 127 && y_pointer == 32)
||(x_pointer == 128 && y_pointer == 32)
||(x_pointer == 129 && y_pointer == 32)
||(x_pointer == 130 && y_pointer == 32)
||(x_pointer == 140 && y_pointer == 32)
||(x_pointer == 141 && y_pointer == 32)
||(x_pointer == 142 && y_pointer == 32)
||(x_pointer == 143 && y_pointer == 32)
||(x_pointer == 144 && y_pointer == 32)
||(x_pointer == 145 && y_pointer == 32)
||(x_pointer == 146 && y_pointer == 32)
||(x_pointer == 147 && y_pointer == 32)
||(x_pointer == 148 && y_pointer == 32)
||(x_pointer == 155 && y_pointer == 32)
||(x_pointer == 156 && y_pointer == 32)
||(x_pointer == 157 && y_pointer == 32)
||(x_pointer == 2 && y_pointer == 33)
||(x_pointer == 3 && y_pointer == 33)
||(x_pointer == 4 && y_pointer == 33)
||(x_pointer == 14 && y_pointer == 33)
||(x_pointer == 15 && y_pointer == 33)
||(x_pointer == 16 && y_pointer == 33)
||(x_pointer == 17 && y_pointer == 33)
||(x_pointer == 18 && y_pointer == 33)
||(x_pointer == 19 && y_pointer == 33)
||(x_pointer == 20 && y_pointer == 33)
||(x_pointer == 21 && y_pointer == 33)
||(x_pointer == 22 && y_pointer == 33)
||(x_pointer == 32 && y_pointer == 33)
||(x_pointer == 33 && y_pointer == 33)
||(x_pointer == 34 && y_pointer == 33)
||(x_pointer == 35 && y_pointer == 33)
||(x_pointer == 36 && y_pointer == 33)
||(x_pointer == 37 && y_pointer == 33)
||(x_pointer == 38 && y_pointer == 33)
||(x_pointer == 39 && y_pointer == 33)
||(x_pointer == 40 && y_pointer == 33)
||(x_pointer == 50 && y_pointer == 33)
||(x_pointer == 51 && y_pointer == 33)
||(x_pointer == 52 && y_pointer == 33)
||(x_pointer == 53 && y_pointer == 33)
||(x_pointer == 54 && y_pointer == 33)
||(x_pointer == 55 && y_pointer == 33)
||(x_pointer == 56 && y_pointer == 33)
||(x_pointer == 57 && y_pointer == 33)
||(x_pointer == 58 && y_pointer == 33)
||(x_pointer == 68 && y_pointer == 33)
||(x_pointer == 69 && y_pointer == 33)
||(x_pointer == 70 && y_pointer == 33)
||(x_pointer == 71 && y_pointer == 33)
||(x_pointer == 72 && y_pointer == 33)
||(x_pointer == 73 && y_pointer == 33)
||(x_pointer == 74 && y_pointer == 33)
||(x_pointer == 75 && y_pointer == 33)
||(x_pointer == 76 && y_pointer == 33)
||(x_pointer == 86 && y_pointer == 33)
||(x_pointer == 87 && y_pointer == 33)
||(x_pointer == 88 && y_pointer == 33)
||(x_pointer == 89 && y_pointer == 33)
||(x_pointer == 90 && y_pointer == 33)
||(x_pointer == 91 && y_pointer == 33)
||(x_pointer == 92 && y_pointer == 33)
||(x_pointer == 93 && y_pointer == 33)
||(x_pointer == 94 && y_pointer == 33)
||(x_pointer == 104 && y_pointer == 33)
||(x_pointer == 105 && y_pointer == 33)
||(x_pointer == 106 && y_pointer == 33)
||(x_pointer == 107 && y_pointer == 33)
||(x_pointer == 108 && y_pointer == 33)
||(x_pointer == 109 && y_pointer == 33)
||(x_pointer == 110 && y_pointer == 33)
||(x_pointer == 111 && y_pointer == 33)
||(x_pointer == 112 && y_pointer == 33)
||(x_pointer == 122 && y_pointer == 33)
||(x_pointer == 123 && y_pointer == 33)
||(x_pointer == 124 && y_pointer == 33)
||(x_pointer == 125 && y_pointer == 33)
||(x_pointer == 126 && y_pointer == 33)
||(x_pointer == 127 && y_pointer == 33)
||(x_pointer == 128 && y_pointer == 33)
||(x_pointer == 129 && y_pointer == 33)
||(x_pointer == 130 && y_pointer == 33)
||(x_pointer == 140 && y_pointer == 33)
||(x_pointer == 141 && y_pointer == 33)
||(x_pointer == 142 && y_pointer == 33)
||(x_pointer == 143 && y_pointer == 33)
||(x_pointer == 144 && y_pointer == 33)
||(x_pointer == 145 && y_pointer == 33)
||(x_pointer == 146 && y_pointer == 33)
||(x_pointer == 147 && y_pointer == 33)
||(x_pointer == 148 && y_pointer == 33)
||(x_pointer == 155 && y_pointer == 33)
||(x_pointer == 156 && y_pointer == 33)
||(x_pointer == 157 && y_pointer == 33)
||(x_pointer == 2 && y_pointer == 34)
||(x_pointer == 3 && y_pointer == 34)
||(x_pointer == 4 && y_pointer == 34)
||(x_pointer == 14 && y_pointer == 34)
||(x_pointer == 15 && y_pointer == 34)
||(x_pointer == 16 && y_pointer == 34)
||(x_pointer == 17 && y_pointer == 34)
||(x_pointer == 18 && y_pointer == 34)
||(x_pointer == 19 && y_pointer == 34)
||(x_pointer == 20 && y_pointer == 34)
||(x_pointer == 21 && y_pointer == 34)
||(x_pointer == 22 && y_pointer == 34)
||(x_pointer == 32 && y_pointer == 34)
||(x_pointer == 33 && y_pointer == 34)
||(x_pointer == 34 && y_pointer == 34)
||(x_pointer == 35 && y_pointer == 34)
||(x_pointer == 36 && y_pointer == 34)
||(x_pointer == 37 && y_pointer == 34)
||(x_pointer == 38 && y_pointer == 34)
||(x_pointer == 39 && y_pointer == 34)
||(x_pointer == 40 && y_pointer == 34)
||(x_pointer == 50 && y_pointer == 34)
||(x_pointer == 51 && y_pointer == 34)
||(x_pointer == 52 && y_pointer == 34)
||(x_pointer == 53 && y_pointer == 34)
||(x_pointer == 54 && y_pointer == 34)
||(x_pointer == 55 && y_pointer == 34)
||(x_pointer == 56 && y_pointer == 34)
||(x_pointer == 57 && y_pointer == 34)
||(x_pointer == 58 && y_pointer == 34)
||(x_pointer == 68 && y_pointer == 34)
||(x_pointer == 69 && y_pointer == 34)
||(x_pointer == 70 && y_pointer == 34)
||(x_pointer == 71 && y_pointer == 34)
||(x_pointer == 72 && y_pointer == 34)
||(x_pointer == 73 && y_pointer == 34)
||(x_pointer == 74 && y_pointer == 34)
||(x_pointer == 75 && y_pointer == 34)
||(x_pointer == 76 && y_pointer == 34)
||(x_pointer == 86 && y_pointer == 34)
||(x_pointer == 87 && y_pointer == 34)
||(x_pointer == 88 && y_pointer == 34)
||(x_pointer == 89 && y_pointer == 34)
||(x_pointer == 90 && y_pointer == 34)
||(x_pointer == 91 && y_pointer == 34)
||(x_pointer == 92 && y_pointer == 34)
||(x_pointer == 93 && y_pointer == 34)
||(x_pointer == 94 && y_pointer == 34)
||(x_pointer == 104 && y_pointer == 34)
||(x_pointer == 105 && y_pointer == 34)
||(x_pointer == 106 && y_pointer == 34)
||(x_pointer == 107 && y_pointer == 34)
||(x_pointer == 108 && y_pointer == 34)
||(x_pointer == 109 && y_pointer == 34)
||(x_pointer == 110 && y_pointer == 34)
||(x_pointer == 111 && y_pointer == 34)
||(x_pointer == 112 && y_pointer == 34)
||(x_pointer == 122 && y_pointer == 34)
||(x_pointer == 123 && y_pointer == 34)
||(x_pointer == 124 && y_pointer == 34)
||(x_pointer == 125 && y_pointer == 34)
||(x_pointer == 126 && y_pointer == 34)
||(x_pointer == 127 && y_pointer == 34)
||(x_pointer == 128 && y_pointer == 34)
||(x_pointer == 129 && y_pointer == 34)
||(x_pointer == 130 && y_pointer == 34)
||(x_pointer == 140 && y_pointer == 34)
||(x_pointer == 141 && y_pointer == 34)
||(x_pointer == 142 && y_pointer == 34)
||(x_pointer == 143 && y_pointer == 34)
||(x_pointer == 144 && y_pointer == 34)
||(x_pointer == 145 && y_pointer == 34)
||(x_pointer == 146 && y_pointer == 34)
||(x_pointer == 147 && y_pointer == 34)
||(x_pointer == 148 && y_pointer == 34)
||(x_pointer == 155 && y_pointer == 34)
||(x_pointer == 156 && y_pointer == 34)
||(x_pointer == 157 && y_pointer == 34)
||(x_pointer == 2 && y_pointer == 35)
||(x_pointer == 3 && y_pointer == 35)
||(x_pointer == 4 && y_pointer == 35)
||(x_pointer == 14 && y_pointer == 35)
||(x_pointer == 15 && y_pointer == 35)
||(x_pointer == 16 && y_pointer == 35)
||(x_pointer == 17 && y_pointer == 35)
||(x_pointer == 18 && y_pointer == 35)
||(x_pointer == 19 && y_pointer == 35)
||(x_pointer == 20 && y_pointer == 35)
||(x_pointer == 21 && y_pointer == 35)
||(x_pointer == 22 && y_pointer == 35)
||(x_pointer == 32 && y_pointer == 35)
||(x_pointer == 33 && y_pointer == 35)
||(x_pointer == 34 && y_pointer == 35)
||(x_pointer == 35 && y_pointer == 35)
||(x_pointer == 36 && y_pointer == 35)
||(x_pointer == 37 && y_pointer == 35)
||(x_pointer == 38 && y_pointer == 35)
||(x_pointer == 39 && y_pointer == 35)
||(x_pointer == 40 && y_pointer == 35)
||(x_pointer == 50 && y_pointer == 35)
||(x_pointer == 51 && y_pointer == 35)
||(x_pointer == 52 && y_pointer == 35)
||(x_pointer == 53 && y_pointer == 35)
||(x_pointer == 54 && y_pointer == 35)
||(x_pointer == 55 && y_pointer == 35)
||(x_pointer == 56 && y_pointer == 35)
||(x_pointer == 57 && y_pointer == 35)
||(x_pointer == 58 && y_pointer == 35)
||(x_pointer == 68 && y_pointer == 35)
||(x_pointer == 69 && y_pointer == 35)
||(x_pointer == 70 && y_pointer == 35)
||(x_pointer == 71 && y_pointer == 35)
||(x_pointer == 72 && y_pointer == 35)
||(x_pointer == 73 && y_pointer == 35)
||(x_pointer == 74 && y_pointer == 35)
||(x_pointer == 75 && y_pointer == 35)
||(x_pointer == 76 && y_pointer == 35)
||(x_pointer == 86 && y_pointer == 35)
||(x_pointer == 87 && y_pointer == 35)
||(x_pointer == 88 && y_pointer == 35)
||(x_pointer == 89 && y_pointer == 35)
||(x_pointer == 90 && y_pointer == 35)
||(x_pointer == 91 && y_pointer == 35)
||(x_pointer == 92 && y_pointer == 35)
||(x_pointer == 93 && y_pointer == 35)
||(x_pointer == 94 && y_pointer == 35)
||(x_pointer == 104 && y_pointer == 35)
||(x_pointer == 105 && y_pointer == 35)
||(x_pointer == 106 && y_pointer == 35)
||(x_pointer == 107 && y_pointer == 35)
||(x_pointer == 108 && y_pointer == 35)
||(x_pointer == 109 && y_pointer == 35)
||(x_pointer == 110 && y_pointer == 35)
||(x_pointer == 111 && y_pointer == 35)
||(x_pointer == 112 && y_pointer == 35)
||(x_pointer == 122 && y_pointer == 35)
||(x_pointer == 123 && y_pointer == 35)
||(x_pointer == 124 && y_pointer == 35)
||(x_pointer == 125 && y_pointer == 35)
||(x_pointer == 126 && y_pointer == 35)
||(x_pointer == 127 && y_pointer == 35)
||(x_pointer == 128 && y_pointer == 35)
||(x_pointer == 129 && y_pointer == 35)
||(x_pointer == 130 && y_pointer == 35)
||(x_pointer == 140 && y_pointer == 35)
||(x_pointer == 141 && y_pointer == 35)
||(x_pointer == 142 && y_pointer == 35)
||(x_pointer == 143 && y_pointer == 35)
||(x_pointer == 144 && y_pointer == 35)
||(x_pointer == 145 && y_pointer == 35)
||(x_pointer == 146 && y_pointer == 35)
||(x_pointer == 147 && y_pointer == 35)
||(x_pointer == 148 && y_pointer == 35)
||(x_pointer == 155 && y_pointer == 35)
||(x_pointer == 156 && y_pointer == 35)
||(x_pointer == 157 && y_pointer == 35)
||(x_pointer == 2 && y_pointer == 36)
||(x_pointer == 3 && y_pointer == 36)
||(x_pointer == 4 && y_pointer == 36)
||(x_pointer == 14 && y_pointer == 36)
||(x_pointer == 15 && y_pointer == 36)
||(x_pointer == 16 && y_pointer == 36)
||(x_pointer == 17 && y_pointer == 36)
||(x_pointer == 18 && y_pointer == 36)
||(x_pointer == 19 && y_pointer == 36)
||(x_pointer == 20 && y_pointer == 36)
||(x_pointer == 21 && y_pointer == 36)
||(x_pointer == 22 && y_pointer == 36)
||(x_pointer == 32 && y_pointer == 36)
||(x_pointer == 33 && y_pointer == 36)
||(x_pointer == 34 && y_pointer == 36)
||(x_pointer == 35 && y_pointer == 36)
||(x_pointer == 36 && y_pointer == 36)
||(x_pointer == 37 && y_pointer == 36)
||(x_pointer == 38 && y_pointer == 36)
||(x_pointer == 39 && y_pointer == 36)
||(x_pointer == 40 && y_pointer == 36)
||(x_pointer == 50 && y_pointer == 36)
||(x_pointer == 51 && y_pointer == 36)
||(x_pointer == 52 && y_pointer == 36)
||(x_pointer == 53 && y_pointer == 36)
||(x_pointer == 54 && y_pointer == 36)
||(x_pointer == 55 && y_pointer == 36)
||(x_pointer == 56 && y_pointer == 36)
||(x_pointer == 57 && y_pointer == 36)
||(x_pointer == 58 && y_pointer == 36)
||(x_pointer == 68 && y_pointer == 36)
||(x_pointer == 69 && y_pointer == 36)
||(x_pointer == 70 && y_pointer == 36)
||(x_pointer == 71 && y_pointer == 36)
||(x_pointer == 72 && y_pointer == 36)
||(x_pointer == 73 && y_pointer == 36)
||(x_pointer == 74 && y_pointer == 36)
||(x_pointer == 75 && y_pointer == 36)
||(x_pointer == 76 && y_pointer == 36)
||(x_pointer == 86 && y_pointer == 36)
||(x_pointer == 87 && y_pointer == 36)
||(x_pointer == 88 && y_pointer == 36)
||(x_pointer == 89 && y_pointer == 36)
||(x_pointer == 90 && y_pointer == 36)
||(x_pointer == 91 && y_pointer == 36)
||(x_pointer == 92 && y_pointer == 36)
||(x_pointer == 93 && y_pointer == 36)
||(x_pointer == 94 && y_pointer == 36)
||(x_pointer == 104 && y_pointer == 36)
||(x_pointer == 105 && y_pointer == 36)
||(x_pointer == 106 && y_pointer == 36)
||(x_pointer == 107 && y_pointer == 36)
||(x_pointer == 108 && y_pointer == 36)
||(x_pointer == 109 && y_pointer == 36)
||(x_pointer == 110 && y_pointer == 36)
||(x_pointer == 111 && y_pointer == 36)
||(x_pointer == 112 && y_pointer == 36)
||(x_pointer == 122 && y_pointer == 36)
||(x_pointer == 123 && y_pointer == 36)
||(x_pointer == 124 && y_pointer == 36)
||(x_pointer == 125 && y_pointer == 36)
||(x_pointer == 126 && y_pointer == 36)
||(x_pointer == 127 && y_pointer == 36)
||(x_pointer == 128 && y_pointer == 36)
||(x_pointer == 129 && y_pointer == 36)
||(x_pointer == 130 && y_pointer == 36)
||(x_pointer == 140 && y_pointer == 36)
||(x_pointer == 141 && y_pointer == 36)
||(x_pointer == 142 && y_pointer == 36)
||(x_pointer == 143 && y_pointer == 36)
||(x_pointer == 144 && y_pointer == 36)
||(x_pointer == 145 && y_pointer == 36)
||(x_pointer == 146 && y_pointer == 36)
||(x_pointer == 147 && y_pointer == 36)
||(x_pointer == 148 && y_pointer == 36)
||(x_pointer == 155 && y_pointer == 36)
||(x_pointer == 156 && y_pointer == 36)
||(x_pointer == 157 && y_pointer == 36)
||(x_pointer == 2 && y_pointer == 37)
||(x_pointer == 3 && y_pointer == 37)
||(x_pointer == 4 && y_pointer == 37)
||(x_pointer == 14 && y_pointer == 37)
||(x_pointer == 15 && y_pointer == 37)
||(x_pointer == 16 && y_pointer == 37)
||(x_pointer == 17 && y_pointer == 37)
||(x_pointer == 18 && y_pointer == 37)
||(x_pointer == 19 && y_pointer == 37)
||(x_pointer == 20 && y_pointer == 37)
||(x_pointer == 21 && y_pointer == 37)
||(x_pointer == 22 && y_pointer == 37)
||(x_pointer == 32 && y_pointer == 37)
||(x_pointer == 33 && y_pointer == 37)
||(x_pointer == 34 && y_pointer == 37)
||(x_pointer == 35 && y_pointer == 37)
||(x_pointer == 36 && y_pointer == 37)
||(x_pointer == 37 && y_pointer == 37)
||(x_pointer == 38 && y_pointer == 37)
||(x_pointer == 39 && y_pointer == 37)
||(x_pointer == 40 && y_pointer == 37)
||(x_pointer == 50 && y_pointer == 37)
||(x_pointer == 51 && y_pointer == 37)
||(x_pointer == 52 && y_pointer == 37)
||(x_pointer == 53 && y_pointer == 37)
||(x_pointer == 54 && y_pointer == 37)
||(x_pointer == 55 && y_pointer == 37)
||(x_pointer == 56 && y_pointer == 37)
||(x_pointer == 57 && y_pointer == 37)
||(x_pointer == 58 && y_pointer == 37)
||(x_pointer == 68 && y_pointer == 37)
||(x_pointer == 69 && y_pointer == 37)
||(x_pointer == 70 && y_pointer == 37)
||(x_pointer == 71 && y_pointer == 37)
||(x_pointer == 72 && y_pointer == 37)
||(x_pointer == 73 && y_pointer == 37)
||(x_pointer == 74 && y_pointer == 37)
||(x_pointer == 75 && y_pointer == 37)
||(x_pointer == 76 && y_pointer == 37)
||(x_pointer == 86 && y_pointer == 37)
||(x_pointer == 87 && y_pointer == 37)
||(x_pointer == 88 && y_pointer == 37)
||(x_pointer == 89 && y_pointer == 37)
||(x_pointer == 90 && y_pointer == 37)
||(x_pointer == 91 && y_pointer == 37)
||(x_pointer == 92 && y_pointer == 37)
||(x_pointer == 93 && y_pointer == 37)
||(x_pointer == 94 && y_pointer == 37)
||(x_pointer == 104 && y_pointer == 37)
||(x_pointer == 105 && y_pointer == 37)
||(x_pointer == 106 && y_pointer == 37)
||(x_pointer == 107 && y_pointer == 37)
||(x_pointer == 108 && y_pointer == 37)
||(x_pointer == 109 && y_pointer == 37)
||(x_pointer == 110 && y_pointer == 37)
||(x_pointer == 111 && y_pointer == 37)
||(x_pointer == 112 && y_pointer == 37)
||(x_pointer == 122 && y_pointer == 37)
||(x_pointer == 123 && y_pointer == 37)
||(x_pointer == 124 && y_pointer == 37)
||(x_pointer == 125 && y_pointer == 37)
||(x_pointer == 126 && y_pointer == 37)
||(x_pointer == 127 && y_pointer == 37)
||(x_pointer == 128 && y_pointer == 37)
||(x_pointer == 129 && y_pointer == 37)
||(x_pointer == 130 && y_pointer == 37)
||(x_pointer == 140 && y_pointer == 37)
||(x_pointer == 141 && y_pointer == 37)
||(x_pointer == 142 && y_pointer == 37)
||(x_pointer == 143 && y_pointer == 37)
||(x_pointer == 144 && y_pointer == 37)
||(x_pointer == 145 && y_pointer == 37)
||(x_pointer == 146 && y_pointer == 37)
||(x_pointer == 147 && y_pointer == 37)
||(x_pointer == 148 && y_pointer == 37)
||(x_pointer == 155 && y_pointer == 37)
||(x_pointer == 156 && y_pointer == 37)
||(x_pointer == 157 && y_pointer == 37)
||(x_pointer == 2 && y_pointer == 38)
||(x_pointer == 3 && y_pointer == 38)
||(x_pointer == 4 && y_pointer == 38)
||(x_pointer == 14 && y_pointer == 38)
||(x_pointer == 15 && y_pointer == 38)
||(x_pointer == 16 && y_pointer == 38)
||(x_pointer == 17 && y_pointer == 38)
||(x_pointer == 18 && y_pointer == 38)
||(x_pointer == 19 && y_pointer == 38)
||(x_pointer == 20 && y_pointer == 38)
||(x_pointer == 21 && y_pointer == 38)
||(x_pointer == 22 && y_pointer == 38)
||(x_pointer == 32 && y_pointer == 38)
||(x_pointer == 33 && y_pointer == 38)
||(x_pointer == 34 && y_pointer == 38)
||(x_pointer == 35 && y_pointer == 38)
||(x_pointer == 36 && y_pointer == 38)
||(x_pointer == 37 && y_pointer == 38)
||(x_pointer == 38 && y_pointer == 38)
||(x_pointer == 39 && y_pointer == 38)
||(x_pointer == 40 && y_pointer == 38)
||(x_pointer == 50 && y_pointer == 38)
||(x_pointer == 51 && y_pointer == 38)
||(x_pointer == 52 && y_pointer == 38)
||(x_pointer == 53 && y_pointer == 38)
||(x_pointer == 54 && y_pointer == 38)
||(x_pointer == 55 && y_pointer == 38)
||(x_pointer == 56 && y_pointer == 38)
||(x_pointer == 57 && y_pointer == 38)
||(x_pointer == 58 && y_pointer == 38)
||(x_pointer == 68 && y_pointer == 38)
||(x_pointer == 69 && y_pointer == 38)
||(x_pointer == 70 && y_pointer == 38)
||(x_pointer == 71 && y_pointer == 38)
||(x_pointer == 72 && y_pointer == 38)
||(x_pointer == 73 && y_pointer == 38)
||(x_pointer == 74 && y_pointer == 38)
||(x_pointer == 75 && y_pointer == 38)
||(x_pointer == 76 && y_pointer == 38)
||(x_pointer == 86 && y_pointer == 38)
||(x_pointer == 87 && y_pointer == 38)
||(x_pointer == 88 && y_pointer == 38)
||(x_pointer == 89 && y_pointer == 38)
||(x_pointer == 90 && y_pointer == 38)
||(x_pointer == 91 && y_pointer == 38)
||(x_pointer == 92 && y_pointer == 38)
||(x_pointer == 93 && y_pointer == 38)
||(x_pointer == 94 && y_pointer == 38)
||(x_pointer == 104 && y_pointer == 38)
||(x_pointer == 105 && y_pointer == 38)
||(x_pointer == 106 && y_pointer == 38)
||(x_pointer == 107 && y_pointer == 38)
||(x_pointer == 108 && y_pointer == 38)
||(x_pointer == 109 && y_pointer == 38)
||(x_pointer == 110 && y_pointer == 38)
||(x_pointer == 111 && y_pointer == 38)
||(x_pointer == 112 && y_pointer == 38)
||(x_pointer == 122 && y_pointer == 38)
||(x_pointer == 123 && y_pointer == 38)
||(x_pointer == 124 && y_pointer == 38)
||(x_pointer == 125 && y_pointer == 38)
||(x_pointer == 126 && y_pointer == 38)
||(x_pointer == 127 && y_pointer == 38)
||(x_pointer == 128 && y_pointer == 38)
||(x_pointer == 129 && y_pointer == 38)
||(x_pointer == 130 && y_pointer == 38)
||(x_pointer == 140 && y_pointer == 38)
||(x_pointer == 141 && y_pointer == 38)
||(x_pointer == 142 && y_pointer == 38)
||(x_pointer == 143 && y_pointer == 38)
||(x_pointer == 144 && y_pointer == 38)
||(x_pointer == 145 && y_pointer == 38)
||(x_pointer == 146 && y_pointer == 38)
||(x_pointer == 147 && y_pointer == 38)
||(x_pointer == 148 && y_pointer == 38)
||(x_pointer == 155 && y_pointer == 38)
||(x_pointer == 156 && y_pointer == 38)
||(x_pointer == 157 && y_pointer == 38)
||(x_pointer == 2 && y_pointer == 39)
||(x_pointer == 3 && y_pointer == 39)
||(x_pointer == 4 && y_pointer == 39)
||(x_pointer == 14 && y_pointer == 39)
||(x_pointer == 15 && y_pointer == 39)
||(x_pointer == 16 && y_pointer == 39)
||(x_pointer == 17 && y_pointer == 39)
||(x_pointer == 18 && y_pointer == 39)
||(x_pointer == 19 && y_pointer == 39)
||(x_pointer == 20 && y_pointer == 39)
||(x_pointer == 21 && y_pointer == 39)
||(x_pointer == 22 && y_pointer == 39)
||(x_pointer == 32 && y_pointer == 39)
||(x_pointer == 33 && y_pointer == 39)
||(x_pointer == 34 && y_pointer == 39)
||(x_pointer == 35 && y_pointer == 39)
||(x_pointer == 36 && y_pointer == 39)
||(x_pointer == 37 && y_pointer == 39)
||(x_pointer == 38 && y_pointer == 39)
||(x_pointer == 39 && y_pointer == 39)
||(x_pointer == 40 && y_pointer == 39)
||(x_pointer == 50 && y_pointer == 39)
||(x_pointer == 51 && y_pointer == 39)
||(x_pointer == 52 && y_pointer == 39)
||(x_pointer == 53 && y_pointer == 39)
||(x_pointer == 54 && y_pointer == 39)
||(x_pointer == 55 && y_pointer == 39)
||(x_pointer == 56 && y_pointer == 39)
||(x_pointer == 57 && y_pointer == 39)
||(x_pointer == 58 && y_pointer == 39)
||(x_pointer == 68 && y_pointer == 39)
||(x_pointer == 69 && y_pointer == 39)
||(x_pointer == 70 && y_pointer == 39)
||(x_pointer == 71 && y_pointer == 39)
||(x_pointer == 72 && y_pointer == 39)
||(x_pointer == 73 && y_pointer == 39)
||(x_pointer == 74 && y_pointer == 39)
||(x_pointer == 75 && y_pointer == 39)
||(x_pointer == 76 && y_pointer == 39)
||(x_pointer == 86 && y_pointer == 39)
||(x_pointer == 87 && y_pointer == 39)
||(x_pointer == 88 && y_pointer == 39)
||(x_pointer == 89 && y_pointer == 39)
||(x_pointer == 90 && y_pointer == 39)
||(x_pointer == 91 && y_pointer == 39)
||(x_pointer == 92 && y_pointer == 39)
||(x_pointer == 93 && y_pointer == 39)
||(x_pointer == 94 && y_pointer == 39)
||(x_pointer == 104 && y_pointer == 39)
||(x_pointer == 105 && y_pointer == 39)
||(x_pointer == 106 && y_pointer == 39)
||(x_pointer == 107 && y_pointer == 39)
||(x_pointer == 108 && y_pointer == 39)
||(x_pointer == 109 && y_pointer == 39)
||(x_pointer == 110 && y_pointer == 39)
||(x_pointer == 111 && y_pointer == 39)
||(x_pointer == 112 && y_pointer == 39)
||(x_pointer == 122 && y_pointer == 39)
||(x_pointer == 123 && y_pointer == 39)
||(x_pointer == 124 && y_pointer == 39)
||(x_pointer == 125 && y_pointer == 39)
||(x_pointer == 126 && y_pointer == 39)
||(x_pointer == 127 && y_pointer == 39)
||(x_pointer == 128 && y_pointer == 39)
||(x_pointer == 129 && y_pointer == 39)
||(x_pointer == 130 && y_pointer == 39)
||(x_pointer == 140 && y_pointer == 39)
||(x_pointer == 141 && y_pointer == 39)
||(x_pointer == 142 && y_pointer == 39)
||(x_pointer == 143 && y_pointer == 39)
||(x_pointer == 144 && y_pointer == 39)
||(x_pointer == 145 && y_pointer == 39)
||(x_pointer == 146 && y_pointer == 39)
||(x_pointer == 147 && y_pointer == 39)
||(x_pointer == 148 && y_pointer == 39)
||(x_pointer == 155 && y_pointer == 39)
||(x_pointer == 156 && y_pointer == 39)
||(x_pointer == 157 && y_pointer == 39)
||(x_pointer == 2 && y_pointer == 40)
||(x_pointer == 3 && y_pointer == 40)
||(x_pointer == 4 && y_pointer == 40)
||(x_pointer == 14 && y_pointer == 40)
||(x_pointer == 15 && y_pointer == 40)
||(x_pointer == 16 && y_pointer == 40)
||(x_pointer == 17 && y_pointer == 40)
||(x_pointer == 18 && y_pointer == 40)
||(x_pointer == 19 && y_pointer == 40)
||(x_pointer == 20 && y_pointer == 40)
||(x_pointer == 21 && y_pointer == 40)
||(x_pointer == 22 && y_pointer == 40)
||(x_pointer == 32 && y_pointer == 40)
||(x_pointer == 33 && y_pointer == 40)
||(x_pointer == 34 && y_pointer == 40)
||(x_pointer == 35 && y_pointer == 40)
||(x_pointer == 36 && y_pointer == 40)
||(x_pointer == 37 && y_pointer == 40)
||(x_pointer == 38 && y_pointer == 40)
||(x_pointer == 39 && y_pointer == 40)
||(x_pointer == 40 && y_pointer == 40)
||(x_pointer == 50 && y_pointer == 40)
||(x_pointer == 51 && y_pointer == 40)
||(x_pointer == 52 && y_pointer == 40)
||(x_pointer == 53 && y_pointer == 40)
||(x_pointer == 54 && y_pointer == 40)
||(x_pointer == 55 && y_pointer == 40)
||(x_pointer == 56 && y_pointer == 40)
||(x_pointer == 57 && y_pointer == 40)
||(x_pointer == 58 && y_pointer == 40)
||(x_pointer == 68 && y_pointer == 40)
||(x_pointer == 69 && y_pointer == 40)
||(x_pointer == 70 && y_pointer == 40)
||(x_pointer == 71 && y_pointer == 40)
||(x_pointer == 72 && y_pointer == 40)
||(x_pointer == 73 && y_pointer == 40)
||(x_pointer == 74 && y_pointer == 40)
||(x_pointer == 75 && y_pointer == 40)
||(x_pointer == 76 && y_pointer == 40)
||(x_pointer == 86 && y_pointer == 40)
||(x_pointer == 87 && y_pointer == 40)
||(x_pointer == 88 && y_pointer == 40)
||(x_pointer == 89 && y_pointer == 40)
||(x_pointer == 90 && y_pointer == 40)
||(x_pointer == 91 && y_pointer == 40)
||(x_pointer == 92 && y_pointer == 40)
||(x_pointer == 93 && y_pointer == 40)
||(x_pointer == 94 && y_pointer == 40)
||(x_pointer == 104 && y_pointer == 40)
||(x_pointer == 105 && y_pointer == 40)
||(x_pointer == 106 && y_pointer == 40)
||(x_pointer == 107 && y_pointer == 40)
||(x_pointer == 108 && y_pointer == 40)
||(x_pointer == 109 && y_pointer == 40)
||(x_pointer == 110 && y_pointer == 40)
||(x_pointer == 111 && y_pointer == 40)
||(x_pointer == 112 && y_pointer == 40)
||(x_pointer == 122 && y_pointer == 40)
||(x_pointer == 123 && y_pointer == 40)
||(x_pointer == 124 && y_pointer == 40)
||(x_pointer == 125 && y_pointer == 40)
||(x_pointer == 126 && y_pointer == 40)
||(x_pointer == 127 && y_pointer == 40)
||(x_pointer == 128 && y_pointer == 40)
||(x_pointer == 129 && y_pointer == 40)
||(x_pointer == 130 && y_pointer == 40)
||(x_pointer == 140 && y_pointer == 40)
||(x_pointer == 141 && y_pointer == 40)
||(x_pointer == 142 && y_pointer == 40)
||(x_pointer == 143 && y_pointer == 40)
||(x_pointer == 144 && y_pointer == 40)
||(x_pointer == 145 && y_pointer == 40)
||(x_pointer == 146 && y_pointer == 40)
||(x_pointer == 147 && y_pointer == 40)
||(x_pointer == 148 && y_pointer == 40)
||(x_pointer == 155 && y_pointer == 40)
||(x_pointer == 156 && y_pointer == 40)
||(x_pointer == 157 && y_pointer == 40)
||(x_pointer == 2 && y_pointer == 41)
||(x_pointer == 3 && y_pointer == 41)
||(x_pointer == 4 && y_pointer == 41)
||(x_pointer == 155 && y_pointer == 41)
||(x_pointer == 156 && y_pointer == 41)
||(x_pointer == 157 && y_pointer == 41)
||(x_pointer == 2 && y_pointer == 42)
||(x_pointer == 3 && y_pointer == 42)
||(x_pointer == 4 && y_pointer == 42)
||(x_pointer == 155 && y_pointer == 42)
||(x_pointer == 156 && y_pointer == 42)
||(x_pointer == 157 && y_pointer == 42)
||(x_pointer == 2 && y_pointer == 43)
||(x_pointer == 3 && y_pointer == 43)
||(x_pointer == 4 && y_pointer == 43)
||(x_pointer == 155 && y_pointer == 43)
||(x_pointer == 156 && y_pointer == 43)
||(x_pointer == 157 && y_pointer == 43)
||(x_pointer == 2 && y_pointer == 44)
||(x_pointer == 3 && y_pointer == 44)
||(x_pointer == 4 && y_pointer == 44)
||(x_pointer == 155 && y_pointer == 44)
||(x_pointer == 156 && y_pointer == 44)
||(x_pointer == 157 && y_pointer == 44)
||(x_pointer == 2 && y_pointer == 45)
||(x_pointer == 3 && y_pointer == 45)
||(x_pointer == 4 && y_pointer == 45)
||(x_pointer == 155 && y_pointer == 45)
||(x_pointer == 156 && y_pointer == 45)
||(x_pointer == 157 && y_pointer == 45)
||(x_pointer == 2 && y_pointer == 46)
||(x_pointer == 3 && y_pointer == 46)
||(x_pointer == 4 && y_pointer == 46)
||(x_pointer == 155 && y_pointer == 46)
||(x_pointer == 156 && y_pointer == 46)
||(x_pointer == 157 && y_pointer == 46)
||(x_pointer == 2 && y_pointer == 47)
||(x_pointer == 3 && y_pointer == 47)
||(x_pointer == 4 && y_pointer == 47)
||(x_pointer == 155 && y_pointer == 47)
||(x_pointer == 156 && y_pointer == 47)
||(x_pointer == 157 && y_pointer == 47)
||(x_pointer == 2 && y_pointer == 48)
||(x_pointer == 3 && y_pointer == 48)
||(x_pointer == 4 && y_pointer == 48)
||(x_pointer == 155 && y_pointer == 48)
||(x_pointer == 156 && y_pointer == 48)
||(x_pointer == 157 && y_pointer == 48)
||(x_pointer == 2 && y_pointer == 49)
||(x_pointer == 3 && y_pointer == 49)
||(x_pointer == 4 && y_pointer == 49)
||(x_pointer == 155 && y_pointer == 49)
||(x_pointer == 156 && y_pointer == 49)
||(x_pointer == 157 && y_pointer == 49)
||(x_pointer == 2 && y_pointer == 50)
||(x_pointer == 3 && y_pointer == 50)
||(x_pointer == 4 && y_pointer == 50)
||(x_pointer == 14 && y_pointer == 50)
||(x_pointer == 15 && y_pointer == 50)
||(x_pointer == 16 && y_pointer == 50)
||(x_pointer == 17 && y_pointer == 50)
||(x_pointer == 18 && y_pointer == 50)
||(x_pointer == 19 && y_pointer == 50)
||(x_pointer == 20 && y_pointer == 50)
||(x_pointer == 21 && y_pointer == 50)
||(x_pointer == 22 && y_pointer == 50)
||(x_pointer == 32 && y_pointer == 50)
||(x_pointer == 33 && y_pointer == 50)
||(x_pointer == 34 && y_pointer == 50)
||(x_pointer == 35 && y_pointer == 50)
||(x_pointer == 36 && y_pointer == 50)
||(x_pointer == 37 && y_pointer == 50)
||(x_pointer == 38 && y_pointer == 50)
||(x_pointer == 39 && y_pointer == 50)
||(x_pointer == 40 && y_pointer == 50)
||(x_pointer == 50 && y_pointer == 50)
||(x_pointer == 51 && y_pointer == 50)
||(x_pointer == 52 && y_pointer == 50)
||(x_pointer == 53 && y_pointer == 50)
||(x_pointer == 54 && y_pointer == 50)
||(x_pointer == 55 && y_pointer == 50)
||(x_pointer == 56 && y_pointer == 50)
||(x_pointer == 57 && y_pointer == 50)
||(x_pointer == 58 && y_pointer == 50)
||(x_pointer == 68 && y_pointer == 50)
||(x_pointer == 69 && y_pointer == 50)
||(x_pointer == 70 && y_pointer == 50)
||(x_pointer == 71 && y_pointer == 50)
||(x_pointer == 72 && y_pointer == 50)
||(x_pointer == 73 && y_pointer == 50)
||(x_pointer == 74 && y_pointer == 50)
||(x_pointer == 75 && y_pointer == 50)
||(x_pointer == 76 && y_pointer == 50)
||(x_pointer == 86 && y_pointer == 50)
||(x_pointer == 87 && y_pointer == 50)
||(x_pointer == 88 && y_pointer == 50)
||(x_pointer == 89 && y_pointer == 50)
||(x_pointer == 90 && y_pointer == 50)
||(x_pointer == 91 && y_pointer == 50)
||(x_pointer == 92 && y_pointer == 50)
||(x_pointer == 93 && y_pointer == 50)
||(x_pointer == 94 && y_pointer == 50)
||(x_pointer == 104 && y_pointer == 50)
||(x_pointer == 105 && y_pointer == 50)
||(x_pointer == 106 && y_pointer == 50)
||(x_pointer == 107 && y_pointer == 50)
||(x_pointer == 108 && y_pointer == 50)
||(x_pointer == 109 && y_pointer == 50)
||(x_pointer == 110 && y_pointer == 50)
||(x_pointer == 111 && y_pointer == 50)
||(x_pointer == 112 && y_pointer == 50)
||(x_pointer == 122 && y_pointer == 50)
||(x_pointer == 123 && y_pointer == 50)
||(x_pointer == 124 && y_pointer == 50)
||(x_pointer == 125 && y_pointer == 50)
||(x_pointer == 126 && y_pointer == 50)
||(x_pointer == 127 && y_pointer == 50)
||(x_pointer == 128 && y_pointer == 50)
||(x_pointer == 129 && y_pointer == 50)
||(x_pointer == 130 && y_pointer == 50)
||(x_pointer == 140 && y_pointer == 50)
||(x_pointer == 141 && y_pointer == 50)
||(x_pointer == 142 && y_pointer == 50)
||(x_pointer == 143 && y_pointer == 50)
||(x_pointer == 144 && y_pointer == 50)
||(x_pointer == 145 && y_pointer == 50)
||(x_pointer == 146 && y_pointer == 50)
||(x_pointer == 147 && y_pointer == 50)
||(x_pointer == 148 && y_pointer == 50)
||(x_pointer == 155 && y_pointer == 50)
||(x_pointer == 156 && y_pointer == 50)
||(x_pointer == 157 && y_pointer == 50)
||(x_pointer == 2 && y_pointer == 51)
||(x_pointer == 3 && y_pointer == 51)
||(x_pointer == 4 && y_pointer == 51)
||(x_pointer == 14 && y_pointer == 51)
||(x_pointer == 15 && y_pointer == 51)
||(x_pointer == 16 && y_pointer == 51)
||(x_pointer == 17 && y_pointer == 51)
||(x_pointer == 18 && y_pointer == 51)
||(x_pointer == 19 && y_pointer == 51)
||(x_pointer == 20 && y_pointer == 51)
||(x_pointer == 21 && y_pointer == 51)
||(x_pointer == 22 && y_pointer == 51)
||(x_pointer == 32 && y_pointer == 51)
||(x_pointer == 33 && y_pointer == 51)
||(x_pointer == 34 && y_pointer == 51)
||(x_pointer == 35 && y_pointer == 51)
||(x_pointer == 36 && y_pointer == 51)
||(x_pointer == 37 && y_pointer == 51)
||(x_pointer == 38 && y_pointer == 51)
||(x_pointer == 39 && y_pointer == 51)
||(x_pointer == 40 && y_pointer == 51)
||(x_pointer == 50 && y_pointer == 51)
||(x_pointer == 51 && y_pointer == 51)
||(x_pointer == 52 && y_pointer == 51)
||(x_pointer == 53 && y_pointer == 51)
||(x_pointer == 54 && y_pointer == 51)
||(x_pointer == 55 && y_pointer == 51)
||(x_pointer == 56 && y_pointer == 51)
||(x_pointer == 57 && y_pointer == 51)
||(x_pointer == 58 && y_pointer == 51)
||(x_pointer == 68 && y_pointer == 51)
||(x_pointer == 69 && y_pointer == 51)
||(x_pointer == 70 && y_pointer == 51)
||(x_pointer == 71 && y_pointer == 51)
||(x_pointer == 72 && y_pointer == 51)
||(x_pointer == 73 && y_pointer == 51)
||(x_pointer == 74 && y_pointer == 51)
||(x_pointer == 75 && y_pointer == 51)
||(x_pointer == 76 && y_pointer == 51)
||(x_pointer == 86 && y_pointer == 51)
||(x_pointer == 87 && y_pointer == 51)
||(x_pointer == 88 && y_pointer == 51)
||(x_pointer == 89 && y_pointer == 51)
||(x_pointer == 90 && y_pointer == 51)
||(x_pointer == 91 && y_pointer == 51)
||(x_pointer == 92 && y_pointer == 51)
||(x_pointer == 93 && y_pointer == 51)
||(x_pointer == 94 && y_pointer == 51)
||(x_pointer == 104 && y_pointer == 51)
||(x_pointer == 105 && y_pointer == 51)
||(x_pointer == 106 && y_pointer == 51)
||(x_pointer == 107 && y_pointer == 51)
||(x_pointer == 108 && y_pointer == 51)
||(x_pointer == 109 && y_pointer == 51)
||(x_pointer == 110 && y_pointer == 51)
||(x_pointer == 111 && y_pointer == 51)
||(x_pointer == 112 && y_pointer == 51)
||(x_pointer == 122 && y_pointer == 51)
||(x_pointer == 123 && y_pointer == 51)
||(x_pointer == 124 && y_pointer == 51)
||(x_pointer == 125 && y_pointer == 51)
||(x_pointer == 126 && y_pointer == 51)
||(x_pointer == 127 && y_pointer == 51)
||(x_pointer == 128 && y_pointer == 51)
||(x_pointer == 129 && y_pointer == 51)
||(x_pointer == 130 && y_pointer == 51)
||(x_pointer == 140 && y_pointer == 51)
||(x_pointer == 141 && y_pointer == 51)
||(x_pointer == 142 && y_pointer == 51)
||(x_pointer == 143 && y_pointer == 51)
||(x_pointer == 144 && y_pointer == 51)
||(x_pointer == 145 && y_pointer == 51)
||(x_pointer == 146 && y_pointer == 51)
||(x_pointer == 147 && y_pointer == 51)
||(x_pointer == 148 && y_pointer == 51)
||(x_pointer == 155 && y_pointer == 51)
||(x_pointer == 156 && y_pointer == 51)
||(x_pointer == 157 && y_pointer == 51)
||(x_pointer == 2 && y_pointer == 52)
||(x_pointer == 3 && y_pointer == 52)
||(x_pointer == 4 && y_pointer == 52)
||(x_pointer == 14 && y_pointer == 52)
||(x_pointer == 15 && y_pointer == 52)
||(x_pointer == 16 && y_pointer == 52)
||(x_pointer == 17 && y_pointer == 52)
||(x_pointer == 18 && y_pointer == 52)
||(x_pointer == 19 && y_pointer == 52)
||(x_pointer == 20 && y_pointer == 52)
||(x_pointer == 21 && y_pointer == 52)
||(x_pointer == 22 && y_pointer == 52)
||(x_pointer == 32 && y_pointer == 52)
||(x_pointer == 33 && y_pointer == 52)
||(x_pointer == 34 && y_pointer == 52)
||(x_pointer == 35 && y_pointer == 52)
||(x_pointer == 36 && y_pointer == 52)
||(x_pointer == 37 && y_pointer == 52)
||(x_pointer == 38 && y_pointer == 52)
||(x_pointer == 39 && y_pointer == 52)
||(x_pointer == 40 && y_pointer == 52)
||(x_pointer == 50 && y_pointer == 52)
||(x_pointer == 51 && y_pointer == 52)
||(x_pointer == 52 && y_pointer == 52)
||(x_pointer == 53 && y_pointer == 52)
||(x_pointer == 54 && y_pointer == 52)
||(x_pointer == 55 && y_pointer == 52)
||(x_pointer == 56 && y_pointer == 52)
||(x_pointer == 57 && y_pointer == 52)
||(x_pointer == 58 && y_pointer == 52)
||(x_pointer == 68 && y_pointer == 52)
||(x_pointer == 69 && y_pointer == 52)
||(x_pointer == 70 && y_pointer == 52)
||(x_pointer == 71 && y_pointer == 52)
||(x_pointer == 72 && y_pointer == 52)
||(x_pointer == 73 && y_pointer == 52)
||(x_pointer == 74 && y_pointer == 52)
||(x_pointer == 75 && y_pointer == 52)
||(x_pointer == 76 && y_pointer == 52)
||(x_pointer == 86 && y_pointer == 52)
||(x_pointer == 87 && y_pointer == 52)
||(x_pointer == 88 && y_pointer == 52)
||(x_pointer == 89 && y_pointer == 52)
||(x_pointer == 90 && y_pointer == 52)
||(x_pointer == 91 && y_pointer == 52)
||(x_pointer == 92 && y_pointer == 52)
||(x_pointer == 93 && y_pointer == 52)
||(x_pointer == 94 && y_pointer == 52)
||(x_pointer == 104 && y_pointer == 52)
||(x_pointer == 105 && y_pointer == 52)
||(x_pointer == 106 && y_pointer == 52)
||(x_pointer == 107 && y_pointer == 52)
||(x_pointer == 108 && y_pointer == 52)
||(x_pointer == 109 && y_pointer == 52)
||(x_pointer == 110 && y_pointer == 52)
||(x_pointer == 111 && y_pointer == 52)
||(x_pointer == 112 && y_pointer == 52)
||(x_pointer == 122 && y_pointer == 52)
||(x_pointer == 123 && y_pointer == 52)
||(x_pointer == 124 && y_pointer == 52)
||(x_pointer == 125 && y_pointer == 52)
||(x_pointer == 126 && y_pointer == 52)
||(x_pointer == 127 && y_pointer == 52)
||(x_pointer == 128 && y_pointer == 52)
||(x_pointer == 129 && y_pointer == 52)
||(x_pointer == 130 && y_pointer == 52)
||(x_pointer == 140 && y_pointer == 52)
||(x_pointer == 141 && y_pointer == 52)
||(x_pointer == 142 && y_pointer == 52)
||(x_pointer == 143 && y_pointer == 52)
||(x_pointer == 144 && y_pointer == 52)
||(x_pointer == 145 && y_pointer == 52)
||(x_pointer == 146 && y_pointer == 52)
||(x_pointer == 147 && y_pointer == 52)
||(x_pointer == 148 && y_pointer == 52)
||(x_pointer == 155 && y_pointer == 52)
||(x_pointer == 156 && y_pointer == 52)
||(x_pointer == 157 && y_pointer == 52)
||(x_pointer == 2 && y_pointer == 53)
||(x_pointer == 3 && y_pointer == 53)
||(x_pointer == 4 && y_pointer == 53)
||(x_pointer == 14 && y_pointer == 53)
||(x_pointer == 15 && y_pointer == 53)
||(x_pointer == 16 && y_pointer == 53)
||(x_pointer == 17 && y_pointer == 53)
||(x_pointer == 18 && y_pointer == 53)
||(x_pointer == 19 && y_pointer == 53)
||(x_pointer == 20 && y_pointer == 53)
||(x_pointer == 21 && y_pointer == 53)
||(x_pointer == 22 && y_pointer == 53)
||(x_pointer == 32 && y_pointer == 53)
||(x_pointer == 33 && y_pointer == 53)
||(x_pointer == 34 && y_pointer == 53)
||(x_pointer == 35 && y_pointer == 53)
||(x_pointer == 36 && y_pointer == 53)
||(x_pointer == 37 && y_pointer == 53)
||(x_pointer == 38 && y_pointer == 53)
||(x_pointer == 39 && y_pointer == 53)
||(x_pointer == 40 && y_pointer == 53)
||(x_pointer == 50 && y_pointer == 53)
||(x_pointer == 51 && y_pointer == 53)
||(x_pointer == 52 && y_pointer == 53)
||(x_pointer == 53 && y_pointer == 53)
||(x_pointer == 54 && y_pointer == 53)
||(x_pointer == 55 && y_pointer == 53)
||(x_pointer == 56 && y_pointer == 53)
||(x_pointer == 57 && y_pointer == 53)
||(x_pointer == 58 && y_pointer == 53)
||(x_pointer == 68 && y_pointer == 53)
||(x_pointer == 69 && y_pointer == 53)
||(x_pointer == 70 && y_pointer == 53)
||(x_pointer == 71 && y_pointer == 53)
||(x_pointer == 72 && y_pointer == 53)
||(x_pointer == 73 && y_pointer == 53)
||(x_pointer == 74 && y_pointer == 53)
||(x_pointer == 75 && y_pointer == 53)
||(x_pointer == 76 && y_pointer == 53)
||(x_pointer == 86 && y_pointer == 53)
||(x_pointer == 87 && y_pointer == 53)
||(x_pointer == 88 && y_pointer == 53)
||(x_pointer == 89 && y_pointer == 53)
||(x_pointer == 90 && y_pointer == 53)
||(x_pointer == 91 && y_pointer == 53)
||(x_pointer == 92 && y_pointer == 53)
||(x_pointer == 93 && y_pointer == 53)
||(x_pointer == 94 && y_pointer == 53)
||(x_pointer == 104 && y_pointer == 53)
||(x_pointer == 105 && y_pointer == 53)
||(x_pointer == 106 && y_pointer == 53)
||(x_pointer == 107 && y_pointer == 53)
||(x_pointer == 108 && y_pointer == 53)
||(x_pointer == 109 && y_pointer == 53)
||(x_pointer == 110 && y_pointer == 53)
||(x_pointer == 111 && y_pointer == 53)
||(x_pointer == 112 && y_pointer == 53)
||(x_pointer == 122 && y_pointer == 53)
||(x_pointer == 123 && y_pointer == 53)
||(x_pointer == 124 && y_pointer == 53)
||(x_pointer == 125 && y_pointer == 53)
||(x_pointer == 126 && y_pointer == 53)
||(x_pointer == 127 && y_pointer == 53)
||(x_pointer == 128 && y_pointer == 53)
||(x_pointer == 129 && y_pointer == 53)
||(x_pointer == 130 && y_pointer == 53)
||(x_pointer == 140 && y_pointer == 53)
||(x_pointer == 141 && y_pointer == 53)
||(x_pointer == 142 && y_pointer == 53)
||(x_pointer == 143 && y_pointer == 53)
||(x_pointer == 144 && y_pointer == 53)
||(x_pointer == 145 && y_pointer == 53)
||(x_pointer == 146 && y_pointer == 53)
||(x_pointer == 147 && y_pointer == 53)
||(x_pointer == 148 && y_pointer == 53)
||(x_pointer == 155 && y_pointer == 53)
||(x_pointer == 156 && y_pointer == 53)
||(x_pointer == 157 && y_pointer == 53)
||(x_pointer == 2 && y_pointer == 54)
||(x_pointer == 3 && y_pointer == 54)
||(x_pointer == 4 && y_pointer == 54)
||(x_pointer == 14 && y_pointer == 54)
||(x_pointer == 15 && y_pointer == 54)
||(x_pointer == 16 && y_pointer == 54)
||(x_pointer == 17 && y_pointer == 54)
||(x_pointer == 18 && y_pointer == 54)
||(x_pointer == 19 && y_pointer == 54)
||(x_pointer == 20 && y_pointer == 54)
||(x_pointer == 21 && y_pointer == 54)
||(x_pointer == 22 && y_pointer == 54)
||(x_pointer == 32 && y_pointer == 54)
||(x_pointer == 33 && y_pointer == 54)
||(x_pointer == 34 && y_pointer == 54)
||(x_pointer == 35 && y_pointer == 54)
||(x_pointer == 36 && y_pointer == 54)
||(x_pointer == 37 && y_pointer == 54)
||(x_pointer == 38 && y_pointer == 54)
||(x_pointer == 39 && y_pointer == 54)
||(x_pointer == 40 && y_pointer == 54)
||(x_pointer == 50 && y_pointer == 54)
||(x_pointer == 51 && y_pointer == 54)
||(x_pointer == 52 && y_pointer == 54)
||(x_pointer == 53 && y_pointer == 54)
||(x_pointer == 54 && y_pointer == 54)
||(x_pointer == 55 && y_pointer == 54)
||(x_pointer == 56 && y_pointer == 54)
||(x_pointer == 57 && y_pointer == 54)
||(x_pointer == 58 && y_pointer == 54)
||(x_pointer == 68 && y_pointer == 54)
||(x_pointer == 69 && y_pointer == 54)
||(x_pointer == 70 && y_pointer == 54)
||(x_pointer == 71 && y_pointer == 54)
||(x_pointer == 72 && y_pointer == 54)
||(x_pointer == 73 && y_pointer == 54)
||(x_pointer == 74 && y_pointer == 54)
||(x_pointer == 75 && y_pointer == 54)
||(x_pointer == 76 && y_pointer == 54)
||(x_pointer == 86 && y_pointer == 54)
||(x_pointer == 87 && y_pointer == 54)
||(x_pointer == 88 && y_pointer == 54)
||(x_pointer == 89 && y_pointer == 54)
||(x_pointer == 90 && y_pointer == 54)
||(x_pointer == 91 && y_pointer == 54)
||(x_pointer == 92 && y_pointer == 54)
||(x_pointer == 93 && y_pointer == 54)
||(x_pointer == 94 && y_pointer == 54)
||(x_pointer == 104 && y_pointer == 54)
||(x_pointer == 105 && y_pointer == 54)
||(x_pointer == 106 && y_pointer == 54)
||(x_pointer == 107 && y_pointer == 54)
||(x_pointer == 108 && y_pointer == 54)
||(x_pointer == 109 && y_pointer == 54)
||(x_pointer == 110 && y_pointer == 54)
||(x_pointer == 111 && y_pointer == 54)
||(x_pointer == 112 && y_pointer == 54)
||(x_pointer == 122 && y_pointer == 54)
||(x_pointer == 123 && y_pointer == 54)
||(x_pointer == 124 && y_pointer == 54)
||(x_pointer == 125 && y_pointer == 54)
||(x_pointer == 126 && y_pointer == 54)
||(x_pointer == 127 && y_pointer == 54)
||(x_pointer == 128 && y_pointer == 54)
||(x_pointer == 129 && y_pointer == 54)
||(x_pointer == 130 && y_pointer == 54)
||(x_pointer == 140 && y_pointer == 54)
||(x_pointer == 141 && y_pointer == 54)
||(x_pointer == 142 && y_pointer == 54)
||(x_pointer == 143 && y_pointer == 54)
||(x_pointer == 144 && y_pointer == 54)
||(x_pointer == 145 && y_pointer == 54)
||(x_pointer == 146 && y_pointer == 54)
||(x_pointer == 147 && y_pointer == 54)
||(x_pointer == 148 && y_pointer == 54)
||(x_pointer == 155 && y_pointer == 54)
||(x_pointer == 156 && y_pointer == 54)
||(x_pointer == 157 && y_pointer == 54)
||(x_pointer == 2 && y_pointer == 55)
||(x_pointer == 3 && y_pointer == 55)
||(x_pointer == 4 && y_pointer == 55)
||(x_pointer == 14 && y_pointer == 55)
||(x_pointer == 15 && y_pointer == 55)
||(x_pointer == 16 && y_pointer == 55)
||(x_pointer == 17 && y_pointer == 55)
||(x_pointer == 18 && y_pointer == 55)
||(x_pointer == 19 && y_pointer == 55)
||(x_pointer == 20 && y_pointer == 55)
||(x_pointer == 21 && y_pointer == 55)
||(x_pointer == 22 && y_pointer == 55)
||(x_pointer == 32 && y_pointer == 55)
||(x_pointer == 33 && y_pointer == 55)
||(x_pointer == 34 && y_pointer == 55)
||(x_pointer == 35 && y_pointer == 55)
||(x_pointer == 36 && y_pointer == 55)
||(x_pointer == 37 && y_pointer == 55)
||(x_pointer == 38 && y_pointer == 55)
||(x_pointer == 39 && y_pointer == 55)
||(x_pointer == 40 && y_pointer == 55)
||(x_pointer == 50 && y_pointer == 55)
||(x_pointer == 51 && y_pointer == 55)
||(x_pointer == 52 && y_pointer == 55)
||(x_pointer == 53 && y_pointer == 55)
||(x_pointer == 54 && y_pointer == 55)
||(x_pointer == 55 && y_pointer == 55)
||(x_pointer == 56 && y_pointer == 55)
||(x_pointer == 57 && y_pointer == 55)
||(x_pointer == 58 && y_pointer == 55)
||(x_pointer == 68 && y_pointer == 55)
||(x_pointer == 69 && y_pointer == 55)
||(x_pointer == 70 && y_pointer == 55)
||(x_pointer == 71 && y_pointer == 55)
||(x_pointer == 72 && y_pointer == 55)
||(x_pointer == 73 && y_pointer == 55)
||(x_pointer == 74 && y_pointer == 55)
||(x_pointer == 75 && y_pointer == 55)
||(x_pointer == 76 && y_pointer == 55)
||(x_pointer == 86 && y_pointer == 55)
||(x_pointer == 87 && y_pointer == 55)
||(x_pointer == 88 && y_pointer == 55)
||(x_pointer == 89 && y_pointer == 55)
||(x_pointer == 90 && y_pointer == 55)
||(x_pointer == 91 && y_pointer == 55)
||(x_pointer == 92 && y_pointer == 55)
||(x_pointer == 93 && y_pointer == 55)
||(x_pointer == 94 && y_pointer == 55)
||(x_pointer == 104 && y_pointer == 55)
||(x_pointer == 105 && y_pointer == 55)
||(x_pointer == 106 && y_pointer == 55)
||(x_pointer == 107 && y_pointer == 55)
||(x_pointer == 108 && y_pointer == 55)
||(x_pointer == 109 && y_pointer == 55)
||(x_pointer == 110 && y_pointer == 55)
||(x_pointer == 111 && y_pointer == 55)
||(x_pointer == 112 && y_pointer == 55)
||(x_pointer == 122 && y_pointer == 55)
||(x_pointer == 123 && y_pointer == 55)
||(x_pointer == 124 && y_pointer == 55)
||(x_pointer == 125 && y_pointer == 55)
||(x_pointer == 126 && y_pointer == 55)
||(x_pointer == 127 && y_pointer == 55)
||(x_pointer == 128 && y_pointer == 55)
||(x_pointer == 129 && y_pointer == 55)
||(x_pointer == 130 && y_pointer == 55)
||(x_pointer == 140 && y_pointer == 55)
||(x_pointer == 141 && y_pointer == 55)
||(x_pointer == 142 && y_pointer == 55)
||(x_pointer == 143 && y_pointer == 55)
||(x_pointer == 144 && y_pointer == 55)
||(x_pointer == 145 && y_pointer == 55)
||(x_pointer == 146 && y_pointer == 55)
||(x_pointer == 147 && y_pointer == 55)
||(x_pointer == 148 && y_pointer == 55)
||(x_pointer == 155 && y_pointer == 55)
||(x_pointer == 156 && y_pointer == 55)
||(x_pointer == 157 && y_pointer == 55)
||(x_pointer == 2 && y_pointer == 56)
||(x_pointer == 3 && y_pointer == 56)
||(x_pointer == 4 && y_pointer == 56)
||(x_pointer == 14 && y_pointer == 56)
||(x_pointer == 15 && y_pointer == 56)
||(x_pointer == 16 && y_pointer == 56)
||(x_pointer == 17 && y_pointer == 56)
||(x_pointer == 18 && y_pointer == 56)
||(x_pointer == 19 && y_pointer == 56)
||(x_pointer == 20 && y_pointer == 56)
||(x_pointer == 21 && y_pointer == 56)
||(x_pointer == 22 && y_pointer == 56)
||(x_pointer == 32 && y_pointer == 56)
||(x_pointer == 33 && y_pointer == 56)
||(x_pointer == 34 && y_pointer == 56)
||(x_pointer == 35 && y_pointer == 56)
||(x_pointer == 36 && y_pointer == 56)
||(x_pointer == 37 && y_pointer == 56)
||(x_pointer == 38 && y_pointer == 56)
||(x_pointer == 39 && y_pointer == 56)
||(x_pointer == 40 && y_pointer == 56)
||(x_pointer == 50 && y_pointer == 56)
||(x_pointer == 51 && y_pointer == 56)
||(x_pointer == 52 && y_pointer == 56)
||(x_pointer == 53 && y_pointer == 56)
||(x_pointer == 54 && y_pointer == 56)
||(x_pointer == 55 && y_pointer == 56)
||(x_pointer == 56 && y_pointer == 56)
||(x_pointer == 57 && y_pointer == 56)
||(x_pointer == 58 && y_pointer == 56)
||(x_pointer == 68 && y_pointer == 56)
||(x_pointer == 69 && y_pointer == 56)
||(x_pointer == 70 && y_pointer == 56)
||(x_pointer == 71 && y_pointer == 56)
||(x_pointer == 72 && y_pointer == 56)
||(x_pointer == 73 && y_pointer == 56)
||(x_pointer == 74 && y_pointer == 56)
||(x_pointer == 75 && y_pointer == 56)
||(x_pointer == 76 && y_pointer == 56)
||(x_pointer == 86 && y_pointer == 56)
||(x_pointer == 87 && y_pointer == 56)
||(x_pointer == 88 && y_pointer == 56)
||(x_pointer == 89 && y_pointer == 56)
||(x_pointer == 90 && y_pointer == 56)
||(x_pointer == 91 && y_pointer == 56)
||(x_pointer == 92 && y_pointer == 56)
||(x_pointer == 93 && y_pointer == 56)
||(x_pointer == 94 && y_pointer == 56)
||(x_pointer == 104 && y_pointer == 56)
||(x_pointer == 105 && y_pointer == 56)
||(x_pointer == 106 && y_pointer == 56)
||(x_pointer == 107 && y_pointer == 56)
||(x_pointer == 108 && y_pointer == 56)
||(x_pointer == 109 && y_pointer == 56)
||(x_pointer == 110 && y_pointer == 56)
||(x_pointer == 111 && y_pointer == 56)
||(x_pointer == 112 && y_pointer == 56)
||(x_pointer == 122 && y_pointer == 56)
||(x_pointer == 123 && y_pointer == 56)
||(x_pointer == 124 && y_pointer == 56)
||(x_pointer == 125 && y_pointer == 56)
||(x_pointer == 126 && y_pointer == 56)
||(x_pointer == 127 && y_pointer == 56)
||(x_pointer == 128 && y_pointer == 56)
||(x_pointer == 129 && y_pointer == 56)
||(x_pointer == 130 && y_pointer == 56)
||(x_pointer == 140 && y_pointer == 56)
||(x_pointer == 141 && y_pointer == 56)
||(x_pointer == 142 && y_pointer == 56)
||(x_pointer == 143 && y_pointer == 56)
||(x_pointer == 144 && y_pointer == 56)
||(x_pointer == 145 && y_pointer == 56)
||(x_pointer == 146 && y_pointer == 56)
||(x_pointer == 147 && y_pointer == 56)
||(x_pointer == 148 && y_pointer == 56)
||(x_pointer == 155 && y_pointer == 56)
||(x_pointer == 156 && y_pointer == 56)
||(x_pointer == 157 && y_pointer == 56)
||(x_pointer == 2 && y_pointer == 57)
||(x_pointer == 3 && y_pointer == 57)
||(x_pointer == 4 && y_pointer == 57)
||(x_pointer == 14 && y_pointer == 57)
||(x_pointer == 15 && y_pointer == 57)
||(x_pointer == 16 && y_pointer == 57)
||(x_pointer == 17 && y_pointer == 57)
||(x_pointer == 18 && y_pointer == 57)
||(x_pointer == 19 && y_pointer == 57)
||(x_pointer == 20 && y_pointer == 57)
||(x_pointer == 21 && y_pointer == 57)
||(x_pointer == 22 && y_pointer == 57)
||(x_pointer == 32 && y_pointer == 57)
||(x_pointer == 33 && y_pointer == 57)
||(x_pointer == 34 && y_pointer == 57)
||(x_pointer == 35 && y_pointer == 57)
||(x_pointer == 36 && y_pointer == 57)
||(x_pointer == 37 && y_pointer == 57)
||(x_pointer == 38 && y_pointer == 57)
||(x_pointer == 39 && y_pointer == 57)
||(x_pointer == 40 && y_pointer == 57)
||(x_pointer == 50 && y_pointer == 57)
||(x_pointer == 51 && y_pointer == 57)
||(x_pointer == 52 && y_pointer == 57)
||(x_pointer == 53 && y_pointer == 57)
||(x_pointer == 54 && y_pointer == 57)
||(x_pointer == 55 && y_pointer == 57)
||(x_pointer == 56 && y_pointer == 57)
||(x_pointer == 57 && y_pointer == 57)
||(x_pointer == 58 && y_pointer == 57)
||(x_pointer == 68 && y_pointer == 57)
||(x_pointer == 69 && y_pointer == 57)
||(x_pointer == 70 && y_pointer == 57)
||(x_pointer == 71 && y_pointer == 57)
||(x_pointer == 72 && y_pointer == 57)
||(x_pointer == 73 && y_pointer == 57)
||(x_pointer == 74 && y_pointer == 57)
||(x_pointer == 75 && y_pointer == 57)
||(x_pointer == 76 && y_pointer == 57)
||(x_pointer == 86 && y_pointer == 57)
||(x_pointer == 87 && y_pointer == 57)
||(x_pointer == 88 && y_pointer == 57)
||(x_pointer == 89 && y_pointer == 57)
||(x_pointer == 90 && y_pointer == 57)
||(x_pointer == 91 && y_pointer == 57)
||(x_pointer == 92 && y_pointer == 57)
||(x_pointer == 93 && y_pointer == 57)
||(x_pointer == 94 && y_pointer == 57)
||(x_pointer == 104 && y_pointer == 57)
||(x_pointer == 105 && y_pointer == 57)
||(x_pointer == 106 && y_pointer == 57)
||(x_pointer == 107 && y_pointer == 57)
||(x_pointer == 108 && y_pointer == 57)
||(x_pointer == 109 && y_pointer == 57)
||(x_pointer == 110 && y_pointer == 57)
||(x_pointer == 111 && y_pointer == 57)
||(x_pointer == 112 && y_pointer == 57)
||(x_pointer == 122 && y_pointer == 57)
||(x_pointer == 123 && y_pointer == 57)
||(x_pointer == 124 && y_pointer == 57)
||(x_pointer == 125 && y_pointer == 57)
||(x_pointer == 126 && y_pointer == 57)
||(x_pointer == 127 && y_pointer == 57)
||(x_pointer == 128 && y_pointer == 57)
||(x_pointer == 129 && y_pointer == 57)
||(x_pointer == 130 && y_pointer == 57)
||(x_pointer == 140 && y_pointer == 57)
||(x_pointer == 141 && y_pointer == 57)
||(x_pointer == 142 && y_pointer == 57)
||(x_pointer == 143 && y_pointer == 57)
||(x_pointer == 144 && y_pointer == 57)
||(x_pointer == 145 && y_pointer == 57)
||(x_pointer == 146 && y_pointer == 57)
||(x_pointer == 147 && y_pointer == 57)
||(x_pointer == 148 && y_pointer == 57)
||(x_pointer == 155 && y_pointer == 57)
||(x_pointer == 156 && y_pointer == 57)
||(x_pointer == 157 && y_pointer == 57)
||(x_pointer == 2 && y_pointer == 58)
||(x_pointer == 3 && y_pointer == 58)
||(x_pointer == 4 && y_pointer == 58)
||(x_pointer == 14 && y_pointer == 58)
||(x_pointer == 15 && y_pointer == 58)
||(x_pointer == 16 && y_pointer == 58)
||(x_pointer == 17 && y_pointer == 58)
||(x_pointer == 18 && y_pointer == 58)
||(x_pointer == 19 && y_pointer == 58)
||(x_pointer == 20 && y_pointer == 58)
||(x_pointer == 21 && y_pointer == 58)
||(x_pointer == 22 && y_pointer == 58)
||(x_pointer == 32 && y_pointer == 58)
||(x_pointer == 33 && y_pointer == 58)
||(x_pointer == 34 && y_pointer == 58)
||(x_pointer == 35 && y_pointer == 58)
||(x_pointer == 36 && y_pointer == 58)
||(x_pointer == 37 && y_pointer == 58)
||(x_pointer == 38 && y_pointer == 58)
||(x_pointer == 39 && y_pointer == 58)
||(x_pointer == 40 && y_pointer == 58)
||(x_pointer == 50 && y_pointer == 58)
||(x_pointer == 51 && y_pointer == 58)
||(x_pointer == 52 && y_pointer == 58)
||(x_pointer == 53 && y_pointer == 58)
||(x_pointer == 54 && y_pointer == 58)
||(x_pointer == 55 && y_pointer == 58)
||(x_pointer == 56 && y_pointer == 58)
||(x_pointer == 57 && y_pointer == 58)
||(x_pointer == 58 && y_pointer == 58)
||(x_pointer == 68 && y_pointer == 58)
||(x_pointer == 69 && y_pointer == 58)
||(x_pointer == 70 && y_pointer == 58)
||(x_pointer == 71 && y_pointer == 58)
||(x_pointer == 72 && y_pointer == 58)
||(x_pointer == 73 && y_pointer == 58)
||(x_pointer == 74 && y_pointer == 58)
||(x_pointer == 75 && y_pointer == 58)
||(x_pointer == 76 && y_pointer == 58)
||(x_pointer == 86 && y_pointer == 58)
||(x_pointer == 87 && y_pointer == 58)
||(x_pointer == 88 && y_pointer == 58)
||(x_pointer == 89 && y_pointer == 58)
||(x_pointer == 90 && y_pointer == 58)
||(x_pointer == 91 && y_pointer == 58)
||(x_pointer == 92 && y_pointer == 58)
||(x_pointer == 93 && y_pointer == 58)
||(x_pointer == 94 && y_pointer == 58)
||(x_pointer == 104 && y_pointer == 58)
||(x_pointer == 105 && y_pointer == 58)
||(x_pointer == 106 && y_pointer == 58)
||(x_pointer == 107 && y_pointer == 58)
||(x_pointer == 108 && y_pointer == 58)
||(x_pointer == 109 && y_pointer == 58)
||(x_pointer == 110 && y_pointer == 58)
||(x_pointer == 111 && y_pointer == 58)
||(x_pointer == 112 && y_pointer == 58)
||(x_pointer == 122 && y_pointer == 58)
||(x_pointer == 123 && y_pointer == 58)
||(x_pointer == 124 && y_pointer == 58)
||(x_pointer == 125 && y_pointer == 58)
||(x_pointer == 126 && y_pointer == 58)
||(x_pointer == 127 && y_pointer == 58)
||(x_pointer == 128 && y_pointer == 58)
||(x_pointer == 129 && y_pointer == 58)
||(x_pointer == 130 && y_pointer == 58)
||(x_pointer == 140 && y_pointer == 58)
||(x_pointer == 141 && y_pointer == 58)
||(x_pointer == 142 && y_pointer == 58)
||(x_pointer == 143 && y_pointer == 58)
||(x_pointer == 144 && y_pointer == 58)
||(x_pointer == 145 && y_pointer == 58)
||(x_pointer == 146 && y_pointer == 58)
||(x_pointer == 147 && y_pointer == 58)
||(x_pointer == 148 && y_pointer == 58)
||(x_pointer == 155 && y_pointer == 58)
||(x_pointer == 156 && y_pointer == 58)
||(x_pointer == 157 && y_pointer == 58)
||(x_pointer == 2 && y_pointer == 59)
||(x_pointer == 3 && y_pointer == 59)
||(x_pointer == 4 && y_pointer == 59)
||(x_pointer == 155 && y_pointer == 59)
||(x_pointer == 156 && y_pointer == 59)
||(x_pointer == 157 && y_pointer == 59)
||(x_pointer == 2 && y_pointer == 60)
||(x_pointer == 3 && y_pointer == 60)
||(x_pointer == 4 && y_pointer == 60)
||(x_pointer == 155 && y_pointer == 60)
||(x_pointer == 156 && y_pointer == 60)
||(x_pointer == 157 && y_pointer == 60)
||(x_pointer == 2 && y_pointer == 61)
||(x_pointer == 3 && y_pointer == 61)
||(x_pointer == 4 && y_pointer == 61)
||(x_pointer == 155 && y_pointer == 61)
||(x_pointer == 156 && y_pointer == 61)
||(x_pointer == 157 && y_pointer == 61)
||(x_pointer == 2 && y_pointer == 62)
||(x_pointer == 3 && y_pointer == 62)
||(x_pointer == 4 && y_pointer == 62)
||(x_pointer == 155 && y_pointer == 62)
||(x_pointer == 156 && y_pointer == 62)
||(x_pointer == 157 && y_pointer == 62)
||(x_pointer == 2 && y_pointer == 63)
||(x_pointer == 3 && y_pointer == 63)
||(x_pointer == 4 && y_pointer == 63)
||(x_pointer == 155 && y_pointer == 63)
||(x_pointer == 156 && y_pointer == 63)
||(x_pointer == 157 && y_pointer == 63)
||(x_pointer == 2 && y_pointer == 64)
||(x_pointer == 3 && y_pointer == 64)
||(x_pointer == 4 && y_pointer == 64)
||(x_pointer == 155 && y_pointer == 64)
||(x_pointer == 156 && y_pointer == 64)
||(x_pointer == 157 && y_pointer == 64)
||(x_pointer == 2 && y_pointer == 65)
||(x_pointer == 3 && y_pointer == 65)
||(x_pointer == 4 && y_pointer == 65)
||(x_pointer == 155 && y_pointer == 65)
||(x_pointer == 156 && y_pointer == 65)
||(x_pointer == 157 && y_pointer == 65)
||(x_pointer == 2 && y_pointer == 66)
||(x_pointer == 3 && y_pointer == 66)
||(x_pointer == 4 && y_pointer == 66)
||(x_pointer == 155 && y_pointer == 66)
||(x_pointer == 156 && y_pointer == 66)
||(x_pointer == 157 && y_pointer == 66)
||(x_pointer == 2 && y_pointer == 67)
||(x_pointer == 3 && y_pointer == 67)
||(x_pointer == 4 && y_pointer == 67)
||(x_pointer == 155 && y_pointer == 67)
||(x_pointer == 156 && y_pointer == 67)
||(x_pointer == 157 && y_pointer == 67)
||(x_pointer == 2 && y_pointer == 68)
||(x_pointer == 3 && y_pointer == 68)
||(x_pointer == 4 && y_pointer == 68)
||(x_pointer == 14 && y_pointer == 68)
||(x_pointer == 15 && y_pointer == 68)
||(x_pointer == 16 && y_pointer == 68)
||(x_pointer == 17 && y_pointer == 68)
||(x_pointer == 18 && y_pointer == 68)
||(x_pointer == 19 && y_pointer == 68)
||(x_pointer == 20 && y_pointer == 68)
||(x_pointer == 21 && y_pointer == 68)
||(x_pointer == 22 && y_pointer == 68)
||(x_pointer == 32 && y_pointer == 68)
||(x_pointer == 33 && y_pointer == 68)
||(x_pointer == 34 && y_pointer == 68)
||(x_pointer == 35 && y_pointer == 68)
||(x_pointer == 36 && y_pointer == 68)
||(x_pointer == 37 && y_pointer == 68)
||(x_pointer == 38 && y_pointer == 68)
||(x_pointer == 39 && y_pointer == 68)
||(x_pointer == 40 && y_pointer == 68)
||(x_pointer == 50 && y_pointer == 68)
||(x_pointer == 51 && y_pointer == 68)
||(x_pointer == 52 && y_pointer == 68)
||(x_pointer == 53 && y_pointer == 68)
||(x_pointer == 54 && y_pointer == 68)
||(x_pointer == 55 && y_pointer == 68)
||(x_pointer == 56 && y_pointer == 68)
||(x_pointer == 57 && y_pointer == 68)
||(x_pointer == 58 && y_pointer == 68)
||(x_pointer == 68 && y_pointer == 68)
||(x_pointer == 69 && y_pointer == 68)
||(x_pointer == 70 && y_pointer == 68)
||(x_pointer == 71 && y_pointer == 68)
||(x_pointer == 72 && y_pointer == 68)
||(x_pointer == 73 && y_pointer == 68)
||(x_pointer == 74 && y_pointer == 68)
||(x_pointer == 75 && y_pointer == 68)
||(x_pointer == 76 && y_pointer == 68)
||(x_pointer == 86 && y_pointer == 68)
||(x_pointer == 87 && y_pointer == 68)
||(x_pointer == 88 && y_pointer == 68)
||(x_pointer == 89 && y_pointer == 68)
||(x_pointer == 90 && y_pointer == 68)
||(x_pointer == 91 && y_pointer == 68)
||(x_pointer == 92 && y_pointer == 68)
||(x_pointer == 93 && y_pointer == 68)
||(x_pointer == 94 && y_pointer == 68)
||(x_pointer == 104 && y_pointer == 68)
||(x_pointer == 105 && y_pointer == 68)
||(x_pointer == 106 && y_pointer == 68)
||(x_pointer == 107 && y_pointer == 68)
||(x_pointer == 108 && y_pointer == 68)
||(x_pointer == 109 && y_pointer == 68)
||(x_pointer == 110 && y_pointer == 68)
||(x_pointer == 111 && y_pointer == 68)
||(x_pointer == 112 && y_pointer == 68)
||(x_pointer == 122 && y_pointer == 68)
||(x_pointer == 123 && y_pointer == 68)
||(x_pointer == 124 && y_pointer == 68)
||(x_pointer == 125 && y_pointer == 68)
||(x_pointer == 126 && y_pointer == 68)
||(x_pointer == 127 && y_pointer == 68)
||(x_pointer == 128 && y_pointer == 68)
||(x_pointer == 129 && y_pointer == 68)
||(x_pointer == 130 && y_pointer == 68)
||(x_pointer == 140 && y_pointer == 68)
||(x_pointer == 141 && y_pointer == 68)
||(x_pointer == 142 && y_pointer == 68)
||(x_pointer == 143 && y_pointer == 68)
||(x_pointer == 144 && y_pointer == 68)
||(x_pointer == 145 && y_pointer == 68)
||(x_pointer == 146 && y_pointer == 68)
||(x_pointer == 147 && y_pointer == 68)
||(x_pointer == 148 && y_pointer == 68)
||(x_pointer == 155 && y_pointer == 68)
||(x_pointer == 156 && y_pointer == 68)
||(x_pointer == 157 && y_pointer == 68)
||(x_pointer == 2 && y_pointer == 69)
||(x_pointer == 3 && y_pointer == 69)
||(x_pointer == 4 && y_pointer == 69)
||(x_pointer == 14 && y_pointer == 69)
||(x_pointer == 15 && y_pointer == 69)
||(x_pointer == 16 && y_pointer == 69)
||(x_pointer == 17 && y_pointer == 69)
||(x_pointer == 18 && y_pointer == 69)
||(x_pointer == 19 && y_pointer == 69)
||(x_pointer == 20 && y_pointer == 69)
||(x_pointer == 21 && y_pointer == 69)
||(x_pointer == 22 && y_pointer == 69)
||(x_pointer == 32 && y_pointer == 69)
||(x_pointer == 33 && y_pointer == 69)
||(x_pointer == 34 && y_pointer == 69)
||(x_pointer == 35 && y_pointer == 69)
||(x_pointer == 36 && y_pointer == 69)
||(x_pointer == 37 && y_pointer == 69)
||(x_pointer == 38 && y_pointer == 69)
||(x_pointer == 39 && y_pointer == 69)
||(x_pointer == 40 && y_pointer == 69)
||(x_pointer == 50 && y_pointer == 69)
||(x_pointer == 51 && y_pointer == 69)
||(x_pointer == 52 && y_pointer == 69)
||(x_pointer == 53 && y_pointer == 69)
||(x_pointer == 54 && y_pointer == 69)
||(x_pointer == 55 && y_pointer == 69)
||(x_pointer == 56 && y_pointer == 69)
||(x_pointer == 57 && y_pointer == 69)
||(x_pointer == 58 && y_pointer == 69)
||(x_pointer == 68 && y_pointer == 69)
||(x_pointer == 69 && y_pointer == 69)
||(x_pointer == 70 && y_pointer == 69)
||(x_pointer == 71 && y_pointer == 69)
||(x_pointer == 72 && y_pointer == 69)
||(x_pointer == 73 && y_pointer == 69)
||(x_pointer == 74 && y_pointer == 69)
||(x_pointer == 75 && y_pointer == 69)
||(x_pointer == 76 && y_pointer == 69)
||(x_pointer == 86 && y_pointer == 69)
||(x_pointer == 87 && y_pointer == 69)
||(x_pointer == 88 && y_pointer == 69)
||(x_pointer == 89 && y_pointer == 69)
||(x_pointer == 90 && y_pointer == 69)
||(x_pointer == 91 && y_pointer == 69)
||(x_pointer == 92 && y_pointer == 69)
||(x_pointer == 93 && y_pointer == 69)
||(x_pointer == 94 && y_pointer == 69)
||(x_pointer == 104 && y_pointer == 69)
||(x_pointer == 105 && y_pointer == 69)
||(x_pointer == 106 && y_pointer == 69)
||(x_pointer == 107 && y_pointer == 69)
||(x_pointer == 108 && y_pointer == 69)
||(x_pointer == 109 && y_pointer == 69)
||(x_pointer == 110 && y_pointer == 69)
||(x_pointer == 111 && y_pointer == 69)
||(x_pointer == 112 && y_pointer == 69)
||(x_pointer == 122 && y_pointer == 69)
||(x_pointer == 123 && y_pointer == 69)
||(x_pointer == 124 && y_pointer == 69)
||(x_pointer == 125 && y_pointer == 69)
||(x_pointer == 126 && y_pointer == 69)
||(x_pointer == 127 && y_pointer == 69)
||(x_pointer == 128 && y_pointer == 69)
||(x_pointer == 129 && y_pointer == 69)
||(x_pointer == 130 && y_pointer == 69)
||(x_pointer == 140 && y_pointer == 69)
||(x_pointer == 141 && y_pointer == 69)
||(x_pointer == 142 && y_pointer == 69)
||(x_pointer == 143 && y_pointer == 69)
||(x_pointer == 144 && y_pointer == 69)
||(x_pointer == 145 && y_pointer == 69)
||(x_pointer == 146 && y_pointer == 69)
||(x_pointer == 147 && y_pointer == 69)
||(x_pointer == 148 && y_pointer == 69)
||(x_pointer == 155 && y_pointer == 69)
||(x_pointer == 156 && y_pointer == 69)
||(x_pointer == 157 && y_pointer == 69)
||(x_pointer == 2 && y_pointer == 70)
||(x_pointer == 3 && y_pointer == 70)
||(x_pointer == 4 && y_pointer == 70)
||(x_pointer == 14 && y_pointer == 70)
||(x_pointer == 15 && y_pointer == 70)
||(x_pointer == 16 && y_pointer == 70)
||(x_pointer == 17 && y_pointer == 70)
||(x_pointer == 18 && y_pointer == 70)
||(x_pointer == 19 && y_pointer == 70)
||(x_pointer == 20 && y_pointer == 70)
||(x_pointer == 21 && y_pointer == 70)
||(x_pointer == 22 && y_pointer == 70)
||(x_pointer == 32 && y_pointer == 70)
||(x_pointer == 33 && y_pointer == 70)
||(x_pointer == 34 && y_pointer == 70)
||(x_pointer == 35 && y_pointer == 70)
||(x_pointer == 36 && y_pointer == 70)
||(x_pointer == 37 && y_pointer == 70)
||(x_pointer == 38 && y_pointer == 70)
||(x_pointer == 39 && y_pointer == 70)
||(x_pointer == 40 && y_pointer == 70)
||(x_pointer == 50 && y_pointer == 70)
||(x_pointer == 51 && y_pointer == 70)
||(x_pointer == 52 && y_pointer == 70)
||(x_pointer == 53 && y_pointer == 70)
||(x_pointer == 54 && y_pointer == 70)
||(x_pointer == 55 && y_pointer == 70)
||(x_pointer == 56 && y_pointer == 70)
||(x_pointer == 57 && y_pointer == 70)
||(x_pointer == 58 && y_pointer == 70)
||(x_pointer == 68 && y_pointer == 70)
||(x_pointer == 69 && y_pointer == 70)
||(x_pointer == 70 && y_pointer == 70)
||(x_pointer == 71 && y_pointer == 70)
||(x_pointer == 72 && y_pointer == 70)
||(x_pointer == 73 && y_pointer == 70)
||(x_pointer == 74 && y_pointer == 70)
||(x_pointer == 75 && y_pointer == 70)
||(x_pointer == 76 && y_pointer == 70)
||(x_pointer == 86 && y_pointer == 70)
||(x_pointer == 87 && y_pointer == 70)
||(x_pointer == 88 && y_pointer == 70)
||(x_pointer == 89 && y_pointer == 70)
||(x_pointer == 90 && y_pointer == 70)
||(x_pointer == 91 && y_pointer == 70)
||(x_pointer == 92 && y_pointer == 70)
||(x_pointer == 93 && y_pointer == 70)
||(x_pointer == 94 && y_pointer == 70)
||(x_pointer == 104 && y_pointer == 70)
||(x_pointer == 105 && y_pointer == 70)
||(x_pointer == 106 && y_pointer == 70)
||(x_pointer == 107 && y_pointer == 70)
||(x_pointer == 108 && y_pointer == 70)
||(x_pointer == 109 && y_pointer == 70)
||(x_pointer == 110 && y_pointer == 70)
||(x_pointer == 111 && y_pointer == 70)
||(x_pointer == 112 && y_pointer == 70)
||(x_pointer == 122 && y_pointer == 70)
||(x_pointer == 123 && y_pointer == 70)
||(x_pointer == 124 && y_pointer == 70)
||(x_pointer == 125 && y_pointer == 70)
||(x_pointer == 126 && y_pointer == 70)
||(x_pointer == 127 && y_pointer == 70)
||(x_pointer == 128 && y_pointer == 70)
||(x_pointer == 129 && y_pointer == 70)
||(x_pointer == 130 && y_pointer == 70)
||(x_pointer == 140 && y_pointer == 70)
||(x_pointer == 141 && y_pointer == 70)
||(x_pointer == 142 && y_pointer == 70)
||(x_pointer == 143 && y_pointer == 70)
||(x_pointer == 144 && y_pointer == 70)
||(x_pointer == 145 && y_pointer == 70)
||(x_pointer == 146 && y_pointer == 70)
||(x_pointer == 147 && y_pointer == 70)
||(x_pointer == 148 && y_pointer == 70)
||(x_pointer == 155 && y_pointer == 70)
||(x_pointer == 156 && y_pointer == 70)
||(x_pointer == 157 && y_pointer == 70)
||(x_pointer == 2 && y_pointer == 71)
||(x_pointer == 3 && y_pointer == 71)
||(x_pointer == 4 && y_pointer == 71)
||(x_pointer == 14 && y_pointer == 71)
||(x_pointer == 15 && y_pointer == 71)
||(x_pointer == 16 && y_pointer == 71)
||(x_pointer == 17 && y_pointer == 71)
||(x_pointer == 18 && y_pointer == 71)
||(x_pointer == 19 && y_pointer == 71)
||(x_pointer == 20 && y_pointer == 71)
||(x_pointer == 21 && y_pointer == 71)
||(x_pointer == 22 && y_pointer == 71)
||(x_pointer == 32 && y_pointer == 71)
||(x_pointer == 33 && y_pointer == 71)
||(x_pointer == 34 && y_pointer == 71)
||(x_pointer == 35 && y_pointer == 71)
||(x_pointer == 36 && y_pointer == 71)
||(x_pointer == 37 && y_pointer == 71)
||(x_pointer == 38 && y_pointer == 71)
||(x_pointer == 39 && y_pointer == 71)
||(x_pointer == 40 && y_pointer == 71)
||(x_pointer == 50 && y_pointer == 71)
||(x_pointer == 51 && y_pointer == 71)
||(x_pointer == 52 && y_pointer == 71)
||(x_pointer == 53 && y_pointer == 71)
||(x_pointer == 54 && y_pointer == 71)
||(x_pointer == 55 && y_pointer == 71)
||(x_pointer == 56 && y_pointer == 71)
||(x_pointer == 57 && y_pointer == 71)
||(x_pointer == 58 && y_pointer == 71)
||(x_pointer == 68 && y_pointer == 71)
||(x_pointer == 69 && y_pointer == 71)
||(x_pointer == 70 && y_pointer == 71)
||(x_pointer == 71 && y_pointer == 71)
||(x_pointer == 72 && y_pointer == 71)
||(x_pointer == 73 && y_pointer == 71)
||(x_pointer == 74 && y_pointer == 71)
||(x_pointer == 75 && y_pointer == 71)
||(x_pointer == 76 && y_pointer == 71)
||(x_pointer == 86 && y_pointer == 71)
||(x_pointer == 87 && y_pointer == 71)
||(x_pointer == 88 && y_pointer == 71)
||(x_pointer == 89 && y_pointer == 71)
||(x_pointer == 90 && y_pointer == 71)
||(x_pointer == 91 && y_pointer == 71)
||(x_pointer == 92 && y_pointer == 71)
||(x_pointer == 93 && y_pointer == 71)
||(x_pointer == 94 && y_pointer == 71)
||(x_pointer == 104 && y_pointer == 71)
||(x_pointer == 105 && y_pointer == 71)
||(x_pointer == 106 && y_pointer == 71)
||(x_pointer == 107 && y_pointer == 71)
||(x_pointer == 108 && y_pointer == 71)
||(x_pointer == 109 && y_pointer == 71)
||(x_pointer == 110 && y_pointer == 71)
||(x_pointer == 111 && y_pointer == 71)
||(x_pointer == 112 && y_pointer == 71)
||(x_pointer == 122 && y_pointer == 71)
||(x_pointer == 123 && y_pointer == 71)
||(x_pointer == 124 && y_pointer == 71)
||(x_pointer == 125 && y_pointer == 71)
||(x_pointer == 126 && y_pointer == 71)
||(x_pointer == 127 && y_pointer == 71)
||(x_pointer == 128 && y_pointer == 71)
||(x_pointer == 129 && y_pointer == 71)
||(x_pointer == 130 && y_pointer == 71)
||(x_pointer == 140 && y_pointer == 71)
||(x_pointer == 141 && y_pointer == 71)
||(x_pointer == 142 && y_pointer == 71)
||(x_pointer == 143 && y_pointer == 71)
||(x_pointer == 144 && y_pointer == 71)
||(x_pointer == 145 && y_pointer == 71)
||(x_pointer == 146 && y_pointer == 71)
||(x_pointer == 147 && y_pointer == 71)
||(x_pointer == 148 && y_pointer == 71)
||(x_pointer == 155 && y_pointer == 71)
||(x_pointer == 156 && y_pointer == 71)
||(x_pointer == 157 && y_pointer == 71)
||(x_pointer == 2 && y_pointer == 72)
||(x_pointer == 3 && y_pointer == 72)
||(x_pointer == 4 && y_pointer == 72)
||(x_pointer == 14 && y_pointer == 72)
||(x_pointer == 15 && y_pointer == 72)
||(x_pointer == 16 && y_pointer == 72)
||(x_pointer == 17 && y_pointer == 72)
||(x_pointer == 18 && y_pointer == 72)
||(x_pointer == 19 && y_pointer == 72)
||(x_pointer == 20 && y_pointer == 72)
||(x_pointer == 21 && y_pointer == 72)
||(x_pointer == 22 && y_pointer == 72)
||(x_pointer == 32 && y_pointer == 72)
||(x_pointer == 33 && y_pointer == 72)
||(x_pointer == 34 && y_pointer == 72)
||(x_pointer == 35 && y_pointer == 72)
||(x_pointer == 36 && y_pointer == 72)
||(x_pointer == 37 && y_pointer == 72)
||(x_pointer == 38 && y_pointer == 72)
||(x_pointer == 39 && y_pointer == 72)
||(x_pointer == 40 && y_pointer == 72)
||(x_pointer == 50 && y_pointer == 72)
||(x_pointer == 51 && y_pointer == 72)
||(x_pointer == 52 && y_pointer == 72)
||(x_pointer == 53 && y_pointer == 72)
||(x_pointer == 54 && y_pointer == 72)
||(x_pointer == 55 && y_pointer == 72)
||(x_pointer == 56 && y_pointer == 72)
||(x_pointer == 57 && y_pointer == 72)
||(x_pointer == 58 && y_pointer == 72)
||(x_pointer == 68 && y_pointer == 72)
||(x_pointer == 69 && y_pointer == 72)
||(x_pointer == 70 && y_pointer == 72)
||(x_pointer == 71 && y_pointer == 72)
||(x_pointer == 72 && y_pointer == 72)
||(x_pointer == 73 && y_pointer == 72)
||(x_pointer == 74 && y_pointer == 72)
||(x_pointer == 75 && y_pointer == 72)
||(x_pointer == 76 && y_pointer == 72)
||(x_pointer == 86 && y_pointer == 72)
||(x_pointer == 87 && y_pointer == 72)
||(x_pointer == 88 && y_pointer == 72)
||(x_pointer == 89 && y_pointer == 72)
||(x_pointer == 90 && y_pointer == 72)
||(x_pointer == 91 && y_pointer == 72)
||(x_pointer == 92 && y_pointer == 72)
||(x_pointer == 93 && y_pointer == 72)
||(x_pointer == 94 && y_pointer == 72)
||(x_pointer == 104 && y_pointer == 72)
||(x_pointer == 105 && y_pointer == 72)
||(x_pointer == 106 && y_pointer == 72)
||(x_pointer == 107 && y_pointer == 72)
||(x_pointer == 108 && y_pointer == 72)
||(x_pointer == 109 && y_pointer == 72)
||(x_pointer == 110 && y_pointer == 72)
||(x_pointer == 111 && y_pointer == 72)
||(x_pointer == 112 && y_pointer == 72)
||(x_pointer == 122 && y_pointer == 72)
||(x_pointer == 123 && y_pointer == 72)
||(x_pointer == 124 && y_pointer == 72)
||(x_pointer == 125 && y_pointer == 72)
||(x_pointer == 126 && y_pointer == 72)
||(x_pointer == 127 && y_pointer == 72)
||(x_pointer == 128 && y_pointer == 72)
||(x_pointer == 129 && y_pointer == 72)
||(x_pointer == 130 && y_pointer == 72)
||(x_pointer == 140 && y_pointer == 72)
||(x_pointer == 141 && y_pointer == 72)
||(x_pointer == 142 && y_pointer == 72)
||(x_pointer == 143 && y_pointer == 72)
||(x_pointer == 144 && y_pointer == 72)
||(x_pointer == 145 && y_pointer == 72)
||(x_pointer == 146 && y_pointer == 72)
||(x_pointer == 147 && y_pointer == 72)
||(x_pointer == 148 && y_pointer == 72)
||(x_pointer == 155 && y_pointer == 72)
||(x_pointer == 156 && y_pointer == 72)
||(x_pointer == 157 && y_pointer == 72)
||(x_pointer == 2 && y_pointer == 73)
||(x_pointer == 3 && y_pointer == 73)
||(x_pointer == 4 && y_pointer == 73)
||(x_pointer == 14 && y_pointer == 73)
||(x_pointer == 15 && y_pointer == 73)
||(x_pointer == 16 && y_pointer == 73)
||(x_pointer == 17 && y_pointer == 73)
||(x_pointer == 18 && y_pointer == 73)
||(x_pointer == 19 && y_pointer == 73)
||(x_pointer == 20 && y_pointer == 73)
||(x_pointer == 21 && y_pointer == 73)
||(x_pointer == 22 && y_pointer == 73)
||(x_pointer == 32 && y_pointer == 73)
||(x_pointer == 33 && y_pointer == 73)
||(x_pointer == 34 && y_pointer == 73)
||(x_pointer == 35 && y_pointer == 73)
||(x_pointer == 36 && y_pointer == 73)
||(x_pointer == 37 && y_pointer == 73)
||(x_pointer == 38 && y_pointer == 73)
||(x_pointer == 39 && y_pointer == 73)
||(x_pointer == 40 && y_pointer == 73)
||(x_pointer == 50 && y_pointer == 73)
||(x_pointer == 51 && y_pointer == 73)
||(x_pointer == 52 && y_pointer == 73)
||(x_pointer == 53 && y_pointer == 73)
||(x_pointer == 54 && y_pointer == 73)
||(x_pointer == 55 && y_pointer == 73)
||(x_pointer == 56 && y_pointer == 73)
||(x_pointer == 57 && y_pointer == 73)
||(x_pointer == 58 && y_pointer == 73)
||(x_pointer == 68 && y_pointer == 73)
||(x_pointer == 69 && y_pointer == 73)
||(x_pointer == 70 && y_pointer == 73)
||(x_pointer == 71 && y_pointer == 73)
||(x_pointer == 72 && y_pointer == 73)
||(x_pointer == 73 && y_pointer == 73)
||(x_pointer == 74 && y_pointer == 73)
||(x_pointer == 75 && y_pointer == 73)
||(x_pointer == 76 && y_pointer == 73)
||(x_pointer == 86 && y_pointer == 73)
||(x_pointer == 87 && y_pointer == 73)
||(x_pointer == 88 && y_pointer == 73)
||(x_pointer == 89 && y_pointer == 73)
||(x_pointer == 90 && y_pointer == 73)
||(x_pointer == 91 && y_pointer == 73)
||(x_pointer == 92 && y_pointer == 73)
||(x_pointer == 93 && y_pointer == 73)
||(x_pointer == 94 && y_pointer == 73)
||(x_pointer == 104 && y_pointer == 73)
||(x_pointer == 105 && y_pointer == 73)
||(x_pointer == 106 && y_pointer == 73)
||(x_pointer == 107 && y_pointer == 73)
||(x_pointer == 108 && y_pointer == 73)
||(x_pointer == 109 && y_pointer == 73)
||(x_pointer == 110 && y_pointer == 73)
||(x_pointer == 111 && y_pointer == 73)
||(x_pointer == 112 && y_pointer == 73)
||(x_pointer == 122 && y_pointer == 73)
||(x_pointer == 123 && y_pointer == 73)
||(x_pointer == 124 && y_pointer == 73)
||(x_pointer == 125 && y_pointer == 73)
||(x_pointer == 126 && y_pointer == 73)
||(x_pointer == 127 && y_pointer == 73)
||(x_pointer == 128 && y_pointer == 73)
||(x_pointer == 129 && y_pointer == 73)
||(x_pointer == 130 && y_pointer == 73)
||(x_pointer == 140 && y_pointer == 73)
||(x_pointer == 141 && y_pointer == 73)
||(x_pointer == 142 && y_pointer == 73)
||(x_pointer == 143 && y_pointer == 73)
||(x_pointer == 144 && y_pointer == 73)
||(x_pointer == 145 && y_pointer == 73)
||(x_pointer == 146 && y_pointer == 73)
||(x_pointer == 147 && y_pointer == 73)
||(x_pointer == 148 && y_pointer == 73)
||(x_pointer == 155 && y_pointer == 73)
||(x_pointer == 156 && y_pointer == 73)
||(x_pointer == 157 && y_pointer == 73)
||(x_pointer == 2 && y_pointer == 74)
||(x_pointer == 3 && y_pointer == 74)
||(x_pointer == 4 && y_pointer == 74)
||(x_pointer == 14 && y_pointer == 74)
||(x_pointer == 15 && y_pointer == 74)
||(x_pointer == 16 && y_pointer == 74)
||(x_pointer == 17 && y_pointer == 74)
||(x_pointer == 18 && y_pointer == 74)
||(x_pointer == 19 && y_pointer == 74)
||(x_pointer == 20 && y_pointer == 74)
||(x_pointer == 21 && y_pointer == 74)
||(x_pointer == 22 && y_pointer == 74)
||(x_pointer == 32 && y_pointer == 74)
||(x_pointer == 33 && y_pointer == 74)
||(x_pointer == 34 && y_pointer == 74)
||(x_pointer == 35 && y_pointer == 74)
||(x_pointer == 36 && y_pointer == 74)
||(x_pointer == 37 && y_pointer == 74)
||(x_pointer == 38 && y_pointer == 74)
||(x_pointer == 39 && y_pointer == 74)
||(x_pointer == 40 && y_pointer == 74)
||(x_pointer == 50 && y_pointer == 74)
||(x_pointer == 51 && y_pointer == 74)
||(x_pointer == 52 && y_pointer == 74)
||(x_pointer == 53 && y_pointer == 74)
||(x_pointer == 54 && y_pointer == 74)
||(x_pointer == 55 && y_pointer == 74)
||(x_pointer == 56 && y_pointer == 74)
||(x_pointer == 57 && y_pointer == 74)
||(x_pointer == 58 && y_pointer == 74)
||(x_pointer == 68 && y_pointer == 74)
||(x_pointer == 69 && y_pointer == 74)
||(x_pointer == 70 && y_pointer == 74)
||(x_pointer == 71 && y_pointer == 74)
||(x_pointer == 72 && y_pointer == 74)
||(x_pointer == 73 && y_pointer == 74)
||(x_pointer == 74 && y_pointer == 74)
||(x_pointer == 75 && y_pointer == 74)
||(x_pointer == 76 && y_pointer == 74)
||(x_pointer == 86 && y_pointer == 74)
||(x_pointer == 87 && y_pointer == 74)
||(x_pointer == 88 && y_pointer == 74)
||(x_pointer == 89 && y_pointer == 74)
||(x_pointer == 90 && y_pointer == 74)
||(x_pointer == 91 && y_pointer == 74)
||(x_pointer == 92 && y_pointer == 74)
||(x_pointer == 93 && y_pointer == 74)
||(x_pointer == 94 && y_pointer == 74)
||(x_pointer == 104 && y_pointer == 74)
||(x_pointer == 105 && y_pointer == 74)
||(x_pointer == 106 && y_pointer == 74)
||(x_pointer == 107 && y_pointer == 74)
||(x_pointer == 108 && y_pointer == 74)
||(x_pointer == 109 && y_pointer == 74)
||(x_pointer == 110 && y_pointer == 74)
||(x_pointer == 111 && y_pointer == 74)
||(x_pointer == 112 && y_pointer == 74)
||(x_pointer == 122 && y_pointer == 74)
||(x_pointer == 123 && y_pointer == 74)
||(x_pointer == 124 && y_pointer == 74)
||(x_pointer == 125 && y_pointer == 74)
||(x_pointer == 126 && y_pointer == 74)
||(x_pointer == 127 && y_pointer == 74)
||(x_pointer == 128 && y_pointer == 74)
||(x_pointer == 129 && y_pointer == 74)
||(x_pointer == 130 && y_pointer == 74)
||(x_pointer == 140 && y_pointer == 74)
||(x_pointer == 141 && y_pointer == 74)
||(x_pointer == 142 && y_pointer == 74)
||(x_pointer == 143 && y_pointer == 74)
||(x_pointer == 144 && y_pointer == 74)
||(x_pointer == 145 && y_pointer == 74)
||(x_pointer == 146 && y_pointer == 74)
||(x_pointer == 147 && y_pointer == 74)
||(x_pointer == 148 && y_pointer == 74)
||(x_pointer == 155 && y_pointer == 74)
||(x_pointer == 156 && y_pointer == 74)
||(x_pointer == 157 && y_pointer == 74)
||(x_pointer == 2 && y_pointer == 75)
||(x_pointer == 3 && y_pointer == 75)
||(x_pointer == 4 && y_pointer == 75)
||(x_pointer == 14 && y_pointer == 75)
||(x_pointer == 15 && y_pointer == 75)
||(x_pointer == 16 && y_pointer == 75)
||(x_pointer == 17 && y_pointer == 75)
||(x_pointer == 18 && y_pointer == 75)
||(x_pointer == 19 && y_pointer == 75)
||(x_pointer == 20 && y_pointer == 75)
||(x_pointer == 21 && y_pointer == 75)
||(x_pointer == 22 && y_pointer == 75)
||(x_pointer == 32 && y_pointer == 75)
||(x_pointer == 33 && y_pointer == 75)
||(x_pointer == 34 && y_pointer == 75)
||(x_pointer == 35 && y_pointer == 75)
||(x_pointer == 36 && y_pointer == 75)
||(x_pointer == 37 && y_pointer == 75)
||(x_pointer == 38 && y_pointer == 75)
||(x_pointer == 39 && y_pointer == 75)
||(x_pointer == 40 && y_pointer == 75)
||(x_pointer == 50 && y_pointer == 75)
||(x_pointer == 51 && y_pointer == 75)
||(x_pointer == 52 && y_pointer == 75)
||(x_pointer == 53 && y_pointer == 75)
||(x_pointer == 54 && y_pointer == 75)
||(x_pointer == 55 && y_pointer == 75)
||(x_pointer == 56 && y_pointer == 75)
||(x_pointer == 57 && y_pointer == 75)
||(x_pointer == 58 && y_pointer == 75)
||(x_pointer == 68 && y_pointer == 75)
||(x_pointer == 69 && y_pointer == 75)
||(x_pointer == 70 && y_pointer == 75)
||(x_pointer == 71 && y_pointer == 75)
||(x_pointer == 72 && y_pointer == 75)
||(x_pointer == 73 && y_pointer == 75)
||(x_pointer == 74 && y_pointer == 75)
||(x_pointer == 75 && y_pointer == 75)
||(x_pointer == 76 && y_pointer == 75)
||(x_pointer == 86 && y_pointer == 75)
||(x_pointer == 87 && y_pointer == 75)
||(x_pointer == 88 && y_pointer == 75)
||(x_pointer == 89 && y_pointer == 75)
||(x_pointer == 90 && y_pointer == 75)
||(x_pointer == 91 && y_pointer == 75)
||(x_pointer == 92 && y_pointer == 75)
||(x_pointer == 93 && y_pointer == 75)
||(x_pointer == 94 && y_pointer == 75)
||(x_pointer == 104 && y_pointer == 75)
||(x_pointer == 105 && y_pointer == 75)
||(x_pointer == 106 && y_pointer == 75)
||(x_pointer == 107 && y_pointer == 75)
||(x_pointer == 108 && y_pointer == 75)
||(x_pointer == 109 && y_pointer == 75)
||(x_pointer == 110 && y_pointer == 75)
||(x_pointer == 111 && y_pointer == 75)
||(x_pointer == 112 && y_pointer == 75)
||(x_pointer == 122 && y_pointer == 75)
||(x_pointer == 123 && y_pointer == 75)
||(x_pointer == 124 && y_pointer == 75)
||(x_pointer == 125 && y_pointer == 75)
||(x_pointer == 126 && y_pointer == 75)
||(x_pointer == 127 && y_pointer == 75)
||(x_pointer == 128 && y_pointer == 75)
||(x_pointer == 129 && y_pointer == 75)
||(x_pointer == 130 && y_pointer == 75)
||(x_pointer == 140 && y_pointer == 75)
||(x_pointer == 141 && y_pointer == 75)
||(x_pointer == 142 && y_pointer == 75)
||(x_pointer == 143 && y_pointer == 75)
||(x_pointer == 144 && y_pointer == 75)
||(x_pointer == 145 && y_pointer == 75)
||(x_pointer == 146 && y_pointer == 75)
||(x_pointer == 147 && y_pointer == 75)
||(x_pointer == 148 && y_pointer == 75)
||(x_pointer == 155 && y_pointer == 75)
||(x_pointer == 156 && y_pointer == 75)
||(x_pointer == 157 && y_pointer == 75)
||(x_pointer == 2 && y_pointer == 76)
||(x_pointer == 3 && y_pointer == 76)
||(x_pointer == 4 && y_pointer == 76)
||(x_pointer == 14 && y_pointer == 76)
||(x_pointer == 15 && y_pointer == 76)
||(x_pointer == 16 && y_pointer == 76)
||(x_pointer == 17 && y_pointer == 76)
||(x_pointer == 18 && y_pointer == 76)
||(x_pointer == 19 && y_pointer == 76)
||(x_pointer == 20 && y_pointer == 76)
||(x_pointer == 21 && y_pointer == 76)
||(x_pointer == 22 && y_pointer == 76)
||(x_pointer == 32 && y_pointer == 76)
||(x_pointer == 33 && y_pointer == 76)
||(x_pointer == 34 && y_pointer == 76)
||(x_pointer == 35 && y_pointer == 76)
||(x_pointer == 36 && y_pointer == 76)
||(x_pointer == 37 && y_pointer == 76)
||(x_pointer == 38 && y_pointer == 76)
||(x_pointer == 39 && y_pointer == 76)
||(x_pointer == 40 && y_pointer == 76)
||(x_pointer == 50 && y_pointer == 76)
||(x_pointer == 51 && y_pointer == 76)
||(x_pointer == 52 && y_pointer == 76)
||(x_pointer == 53 && y_pointer == 76)
||(x_pointer == 54 && y_pointer == 76)
||(x_pointer == 55 && y_pointer == 76)
||(x_pointer == 56 && y_pointer == 76)
||(x_pointer == 57 && y_pointer == 76)
||(x_pointer == 58 && y_pointer == 76)
||(x_pointer == 68 && y_pointer == 76)
||(x_pointer == 69 && y_pointer == 76)
||(x_pointer == 70 && y_pointer == 76)
||(x_pointer == 71 && y_pointer == 76)
||(x_pointer == 72 && y_pointer == 76)
||(x_pointer == 73 && y_pointer == 76)
||(x_pointer == 74 && y_pointer == 76)
||(x_pointer == 75 && y_pointer == 76)
||(x_pointer == 76 && y_pointer == 76)
||(x_pointer == 86 && y_pointer == 76)
||(x_pointer == 87 && y_pointer == 76)
||(x_pointer == 88 && y_pointer == 76)
||(x_pointer == 89 && y_pointer == 76)
||(x_pointer == 90 && y_pointer == 76)
||(x_pointer == 91 && y_pointer == 76)
||(x_pointer == 92 && y_pointer == 76)
||(x_pointer == 93 && y_pointer == 76)
||(x_pointer == 94 && y_pointer == 76)
||(x_pointer == 104 && y_pointer == 76)
||(x_pointer == 105 && y_pointer == 76)
||(x_pointer == 106 && y_pointer == 76)
||(x_pointer == 107 && y_pointer == 76)
||(x_pointer == 108 && y_pointer == 76)
||(x_pointer == 109 && y_pointer == 76)
||(x_pointer == 110 && y_pointer == 76)
||(x_pointer == 111 && y_pointer == 76)
||(x_pointer == 112 && y_pointer == 76)
||(x_pointer == 122 && y_pointer == 76)
||(x_pointer == 123 && y_pointer == 76)
||(x_pointer == 124 && y_pointer == 76)
||(x_pointer == 125 && y_pointer == 76)
||(x_pointer == 126 && y_pointer == 76)
||(x_pointer == 127 && y_pointer == 76)
||(x_pointer == 128 && y_pointer == 76)
||(x_pointer == 129 && y_pointer == 76)
||(x_pointer == 130 && y_pointer == 76)
||(x_pointer == 140 && y_pointer == 76)
||(x_pointer == 141 && y_pointer == 76)
||(x_pointer == 142 && y_pointer == 76)
||(x_pointer == 143 && y_pointer == 76)
||(x_pointer == 144 && y_pointer == 76)
||(x_pointer == 145 && y_pointer == 76)
||(x_pointer == 146 && y_pointer == 76)
||(x_pointer == 147 && y_pointer == 76)
||(x_pointer == 148 && y_pointer == 76)
||(x_pointer == 155 && y_pointer == 76)
||(x_pointer == 156 && y_pointer == 76)
||(x_pointer == 157 && y_pointer == 76)
||(x_pointer == 2 && y_pointer == 77)
||(x_pointer == 3 && y_pointer == 77)
||(x_pointer == 4 && y_pointer == 77)
||(x_pointer == 155 && y_pointer == 77)
||(x_pointer == 156 && y_pointer == 77)
||(x_pointer == 157 && y_pointer == 77)
||(x_pointer == 2 && y_pointer == 78)
||(x_pointer == 3 && y_pointer == 78)
||(x_pointer == 4 && y_pointer == 78)
||(x_pointer == 155 && y_pointer == 78)
||(x_pointer == 156 && y_pointer == 78)
||(x_pointer == 157 && y_pointer == 78)
||(x_pointer == 2 && y_pointer == 79)
||(x_pointer == 3 && y_pointer == 79)
||(x_pointer == 4 && y_pointer == 79)
||(x_pointer == 155 && y_pointer == 79)
||(x_pointer == 156 && y_pointer == 79)
||(x_pointer == 157 && y_pointer == 79)
||(x_pointer == 2 && y_pointer == 80)
||(x_pointer == 3 && y_pointer == 80)
||(x_pointer == 4 && y_pointer == 80)
||(x_pointer == 155 && y_pointer == 80)
||(x_pointer == 156 && y_pointer == 80)
||(x_pointer == 157 && y_pointer == 80)
||(x_pointer == 2 && y_pointer == 81)
||(x_pointer == 3 && y_pointer == 81)
||(x_pointer == 4 && y_pointer == 81)
||(x_pointer == 155 && y_pointer == 81)
||(x_pointer == 156 && y_pointer == 81)
||(x_pointer == 157 && y_pointer == 81)
||(x_pointer == 2 && y_pointer == 82)
||(x_pointer == 3 && y_pointer == 82)
||(x_pointer == 4 && y_pointer == 82)
||(x_pointer == 155 && y_pointer == 82)
||(x_pointer == 156 && y_pointer == 82)
||(x_pointer == 157 && y_pointer == 82)
||(x_pointer == 2 && y_pointer == 83)
||(x_pointer == 3 && y_pointer == 83)
||(x_pointer == 4 && y_pointer == 83)
||(x_pointer == 155 && y_pointer == 83)
||(x_pointer == 156 && y_pointer == 83)
||(x_pointer == 157 && y_pointer == 83)
||(x_pointer == 2 && y_pointer == 84)
||(x_pointer == 3 && y_pointer == 84)
||(x_pointer == 4 && y_pointer == 84)
||(x_pointer == 155 && y_pointer == 84)
||(x_pointer == 156 && y_pointer == 84)
||(x_pointer == 157 && y_pointer == 84)
||(x_pointer == 2 && y_pointer == 85)
||(x_pointer == 3 && y_pointer == 85)
||(x_pointer == 4 && y_pointer == 85)
||(x_pointer == 155 && y_pointer == 85)
||(x_pointer == 156 && y_pointer == 85)
||(x_pointer == 157 && y_pointer == 85)
||(x_pointer == 2 && y_pointer == 86)
||(x_pointer == 3 && y_pointer == 86)
||(x_pointer == 4 && y_pointer == 86)
||(x_pointer == 14 && y_pointer == 86)
||(x_pointer == 15 && y_pointer == 86)
||(x_pointer == 16 && y_pointer == 86)
||(x_pointer == 17 && y_pointer == 86)
||(x_pointer == 18 && y_pointer == 86)
||(x_pointer == 19 && y_pointer == 86)
||(x_pointer == 20 && y_pointer == 86)
||(x_pointer == 21 && y_pointer == 86)
||(x_pointer == 22 && y_pointer == 86)
||(x_pointer == 32 && y_pointer == 86)
||(x_pointer == 33 && y_pointer == 86)
||(x_pointer == 34 && y_pointer == 86)
||(x_pointer == 35 && y_pointer == 86)
||(x_pointer == 36 && y_pointer == 86)
||(x_pointer == 37 && y_pointer == 86)
||(x_pointer == 38 && y_pointer == 86)
||(x_pointer == 39 && y_pointer == 86)
||(x_pointer == 40 && y_pointer == 86)
||(x_pointer == 50 && y_pointer == 86)
||(x_pointer == 51 && y_pointer == 86)
||(x_pointer == 52 && y_pointer == 86)
||(x_pointer == 53 && y_pointer == 86)
||(x_pointer == 54 && y_pointer == 86)
||(x_pointer == 55 && y_pointer == 86)
||(x_pointer == 56 && y_pointer == 86)
||(x_pointer == 57 && y_pointer == 86)
||(x_pointer == 58 && y_pointer == 86)
||(x_pointer == 68 && y_pointer == 86)
||(x_pointer == 69 && y_pointer == 86)
||(x_pointer == 70 && y_pointer == 86)
||(x_pointer == 71 && y_pointer == 86)
||(x_pointer == 72 && y_pointer == 86)
||(x_pointer == 73 && y_pointer == 86)
||(x_pointer == 74 && y_pointer == 86)
||(x_pointer == 75 && y_pointer == 86)
||(x_pointer == 76 && y_pointer == 86)
||(x_pointer == 86 && y_pointer == 86)
||(x_pointer == 87 && y_pointer == 86)
||(x_pointer == 88 && y_pointer == 86)
||(x_pointer == 89 && y_pointer == 86)
||(x_pointer == 90 && y_pointer == 86)
||(x_pointer == 91 && y_pointer == 86)
||(x_pointer == 92 && y_pointer == 86)
||(x_pointer == 93 && y_pointer == 86)
||(x_pointer == 94 && y_pointer == 86)
||(x_pointer == 104 && y_pointer == 86)
||(x_pointer == 105 && y_pointer == 86)
||(x_pointer == 106 && y_pointer == 86)
||(x_pointer == 107 && y_pointer == 86)
||(x_pointer == 108 && y_pointer == 86)
||(x_pointer == 109 && y_pointer == 86)
||(x_pointer == 110 && y_pointer == 86)
||(x_pointer == 111 && y_pointer == 86)
||(x_pointer == 112 && y_pointer == 86)
||(x_pointer == 122 && y_pointer == 86)
||(x_pointer == 123 && y_pointer == 86)
||(x_pointer == 124 && y_pointer == 86)
||(x_pointer == 125 && y_pointer == 86)
||(x_pointer == 126 && y_pointer == 86)
||(x_pointer == 127 && y_pointer == 86)
||(x_pointer == 128 && y_pointer == 86)
||(x_pointer == 129 && y_pointer == 86)
||(x_pointer == 130 && y_pointer == 86)
||(x_pointer == 140 && y_pointer == 86)
||(x_pointer == 141 && y_pointer == 86)
||(x_pointer == 142 && y_pointer == 86)
||(x_pointer == 143 && y_pointer == 86)
||(x_pointer == 144 && y_pointer == 86)
||(x_pointer == 145 && y_pointer == 86)
||(x_pointer == 146 && y_pointer == 86)
||(x_pointer == 147 && y_pointer == 86)
||(x_pointer == 148 && y_pointer == 86)
||(x_pointer == 155 && y_pointer == 86)
||(x_pointer == 156 && y_pointer == 86)
||(x_pointer == 157 && y_pointer == 86)
||(x_pointer == 2 && y_pointer == 87)
||(x_pointer == 3 && y_pointer == 87)
||(x_pointer == 4 && y_pointer == 87)
||(x_pointer == 14 && y_pointer == 87)
||(x_pointer == 15 && y_pointer == 87)
||(x_pointer == 16 && y_pointer == 87)
||(x_pointer == 17 && y_pointer == 87)
||(x_pointer == 18 && y_pointer == 87)
||(x_pointer == 19 && y_pointer == 87)
||(x_pointer == 20 && y_pointer == 87)
||(x_pointer == 21 && y_pointer == 87)
||(x_pointer == 22 && y_pointer == 87)
||(x_pointer == 32 && y_pointer == 87)
||(x_pointer == 33 && y_pointer == 87)
||(x_pointer == 34 && y_pointer == 87)
||(x_pointer == 35 && y_pointer == 87)
||(x_pointer == 36 && y_pointer == 87)
||(x_pointer == 37 && y_pointer == 87)
||(x_pointer == 38 && y_pointer == 87)
||(x_pointer == 39 && y_pointer == 87)
||(x_pointer == 40 && y_pointer == 87)
||(x_pointer == 50 && y_pointer == 87)
||(x_pointer == 51 && y_pointer == 87)
||(x_pointer == 52 && y_pointer == 87)
||(x_pointer == 53 && y_pointer == 87)
||(x_pointer == 54 && y_pointer == 87)
||(x_pointer == 55 && y_pointer == 87)
||(x_pointer == 56 && y_pointer == 87)
||(x_pointer == 57 && y_pointer == 87)
||(x_pointer == 58 && y_pointer == 87)
||(x_pointer == 68 && y_pointer == 87)
||(x_pointer == 69 && y_pointer == 87)
||(x_pointer == 70 && y_pointer == 87)
||(x_pointer == 71 && y_pointer == 87)
||(x_pointer == 72 && y_pointer == 87)
||(x_pointer == 73 && y_pointer == 87)
||(x_pointer == 74 && y_pointer == 87)
||(x_pointer == 75 && y_pointer == 87)
||(x_pointer == 76 && y_pointer == 87)
||(x_pointer == 86 && y_pointer == 87)
||(x_pointer == 87 && y_pointer == 87)
||(x_pointer == 88 && y_pointer == 87)
||(x_pointer == 89 && y_pointer == 87)
||(x_pointer == 90 && y_pointer == 87)
||(x_pointer == 91 && y_pointer == 87)
||(x_pointer == 92 && y_pointer == 87)
||(x_pointer == 93 && y_pointer == 87)
||(x_pointer == 94 && y_pointer == 87)
||(x_pointer == 104 && y_pointer == 87)
||(x_pointer == 105 && y_pointer == 87)
||(x_pointer == 106 && y_pointer == 87)
||(x_pointer == 107 && y_pointer == 87)
||(x_pointer == 108 && y_pointer == 87)
||(x_pointer == 109 && y_pointer == 87)
||(x_pointer == 110 && y_pointer == 87)
||(x_pointer == 111 && y_pointer == 87)
||(x_pointer == 112 && y_pointer == 87)
||(x_pointer == 122 && y_pointer == 87)
||(x_pointer == 123 && y_pointer == 87)
||(x_pointer == 124 && y_pointer == 87)
||(x_pointer == 125 && y_pointer == 87)
||(x_pointer == 126 && y_pointer == 87)
||(x_pointer == 127 && y_pointer == 87)
||(x_pointer == 128 && y_pointer == 87)
||(x_pointer == 129 && y_pointer == 87)
||(x_pointer == 130 && y_pointer == 87)
||(x_pointer == 140 && y_pointer == 87)
||(x_pointer == 141 && y_pointer == 87)
||(x_pointer == 142 && y_pointer == 87)
||(x_pointer == 143 && y_pointer == 87)
||(x_pointer == 144 && y_pointer == 87)
||(x_pointer == 145 && y_pointer == 87)
||(x_pointer == 146 && y_pointer == 87)
||(x_pointer == 147 && y_pointer == 87)
||(x_pointer == 148 && y_pointer == 87)
||(x_pointer == 155 && y_pointer == 87)
||(x_pointer == 156 && y_pointer == 87)
||(x_pointer == 157 && y_pointer == 87)
||(x_pointer == 2 && y_pointer == 88)
||(x_pointer == 3 && y_pointer == 88)
||(x_pointer == 4 && y_pointer == 88)
||(x_pointer == 14 && y_pointer == 88)
||(x_pointer == 15 && y_pointer == 88)
||(x_pointer == 16 && y_pointer == 88)
||(x_pointer == 17 && y_pointer == 88)
||(x_pointer == 18 && y_pointer == 88)
||(x_pointer == 19 && y_pointer == 88)
||(x_pointer == 20 && y_pointer == 88)
||(x_pointer == 21 && y_pointer == 88)
||(x_pointer == 22 && y_pointer == 88)
||(x_pointer == 32 && y_pointer == 88)
||(x_pointer == 33 && y_pointer == 88)
||(x_pointer == 34 && y_pointer == 88)
||(x_pointer == 35 && y_pointer == 88)
||(x_pointer == 36 && y_pointer == 88)
||(x_pointer == 37 && y_pointer == 88)
||(x_pointer == 38 && y_pointer == 88)
||(x_pointer == 39 && y_pointer == 88)
||(x_pointer == 40 && y_pointer == 88)
||(x_pointer == 50 && y_pointer == 88)
||(x_pointer == 51 && y_pointer == 88)
||(x_pointer == 52 && y_pointer == 88)
||(x_pointer == 53 && y_pointer == 88)
||(x_pointer == 54 && y_pointer == 88)
||(x_pointer == 55 && y_pointer == 88)
||(x_pointer == 56 && y_pointer == 88)
||(x_pointer == 57 && y_pointer == 88)
||(x_pointer == 58 && y_pointer == 88)
||(x_pointer == 68 && y_pointer == 88)
||(x_pointer == 69 && y_pointer == 88)
||(x_pointer == 70 && y_pointer == 88)
||(x_pointer == 71 && y_pointer == 88)
||(x_pointer == 72 && y_pointer == 88)
||(x_pointer == 73 && y_pointer == 88)
||(x_pointer == 74 && y_pointer == 88)
||(x_pointer == 75 && y_pointer == 88)
||(x_pointer == 76 && y_pointer == 88)
||(x_pointer == 86 && y_pointer == 88)
||(x_pointer == 87 && y_pointer == 88)
||(x_pointer == 88 && y_pointer == 88)
||(x_pointer == 89 && y_pointer == 88)
||(x_pointer == 90 && y_pointer == 88)
||(x_pointer == 91 && y_pointer == 88)
||(x_pointer == 92 && y_pointer == 88)
||(x_pointer == 93 && y_pointer == 88)
||(x_pointer == 94 && y_pointer == 88)
||(x_pointer == 104 && y_pointer == 88)
||(x_pointer == 105 && y_pointer == 88)
||(x_pointer == 106 && y_pointer == 88)
||(x_pointer == 107 && y_pointer == 88)
||(x_pointer == 108 && y_pointer == 88)
||(x_pointer == 109 && y_pointer == 88)
||(x_pointer == 110 && y_pointer == 88)
||(x_pointer == 111 && y_pointer == 88)
||(x_pointer == 112 && y_pointer == 88)
||(x_pointer == 122 && y_pointer == 88)
||(x_pointer == 123 && y_pointer == 88)
||(x_pointer == 124 && y_pointer == 88)
||(x_pointer == 125 && y_pointer == 88)
||(x_pointer == 126 && y_pointer == 88)
||(x_pointer == 127 && y_pointer == 88)
||(x_pointer == 128 && y_pointer == 88)
||(x_pointer == 129 && y_pointer == 88)
||(x_pointer == 130 && y_pointer == 88)
||(x_pointer == 140 && y_pointer == 88)
||(x_pointer == 141 && y_pointer == 88)
||(x_pointer == 142 && y_pointer == 88)
||(x_pointer == 143 && y_pointer == 88)
||(x_pointer == 144 && y_pointer == 88)
||(x_pointer == 145 && y_pointer == 88)
||(x_pointer == 146 && y_pointer == 88)
||(x_pointer == 147 && y_pointer == 88)
||(x_pointer == 148 && y_pointer == 88)
||(x_pointer == 155 && y_pointer == 88)
||(x_pointer == 156 && y_pointer == 88)
||(x_pointer == 157 && y_pointer == 88)
||(x_pointer == 2 && y_pointer == 89)
||(x_pointer == 3 && y_pointer == 89)
||(x_pointer == 4 && y_pointer == 89)
||(x_pointer == 14 && y_pointer == 89)
||(x_pointer == 15 && y_pointer == 89)
||(x_pointer == 16 && y_pointer == 89)
||(x_pointer == 17 && y_pointer == 89)
||(x_pointer == 18 && y_pointer == 89)
||(x_pointer == 19 && y_pointer == 89)
||(x_pointer == 20 && y_pointer == 89)
||(x_pointer == 21 && y_pointer == 89)
||(x_pointer == 22 && y_pointer == 89)
||(x_pointer == 32 && y_pointer == 89)
||(x_pointer == 33 && y_pointer == 89)
||(x_pointer == 34 && y_pointer == 89)
||(x_pointer == 35 && y_pointer == 89)
||(x_pointer == 36 && y_pointer == 89)
||(x_pointer == 37 && y_pointer == 89)
||(x_pointer == 38 && y_pointer == 89)
||(x_pointer == 39 && y_pointer == 89)
||(x_pointer == 40 && y_pointer == 89)
||(x_pointer == 50 && y_pointer == 89)
||(x_pointer == 51 && y_pointer == 89)
||(x_pointer == 52 && y_pointer == 89)
||(x_pointer == 53 && y_pointer == 89)
||(x_pointer == 54 && y_pointer == 89)
||(x_pointer == 55 && y_pointer == 89)
||(x_pointer == 56 && y_pointer == 89)
||(x_pointer == 57 && y_pointer == 89)
||(x_pointer == 58 && y_pointer == 89)
||(x_pointer == 68 && y_pointer == 89)
||(x_pointer == 69 && y_pointer == 89)
||(x_pointer == 70 && y_pointer == 89)
||(x_pointer == 71 && y_pointer == 89)
||(x_pointer == 72 && y_pointer == 89)
||(x_pointer == 73 && y_pointer == 89)
||(x_pointer == 74 && y_pointer == 89)
||(x_pointer == 75 && y_pointer == 89)
||(x_pointer == 76 && y_pointer == 89)
||(x_pointer == 86 && y_pointer == 89)
||(x_pointer == 87 && y_pointer == 89)
||(x_pointer == 88 && y_pointer == 89)
||(x_pointer == 89 && y_pointer == 89)
||(x_pointer == 90 && y_pointer == 89)
||(x_pointer == 91 && y_pointer == 89)
||(x_pointer == 92 && y_pointer == 89)
||(x_pointer == 93 && y_pointer == 89)
||(x_pointer == 94 && y_pointer == 89)
||(x_pointer == 104 && y_pointer == 89)
||(x_pointer == 105 && y_pointer == 89)
||(x_pointer == 106 && y_pointer == 89)
||(x_pointer == 107 && y_pointer == 89)
||(x_pointer == 108 && y_pointer == 89)
||(x_pointer == 109 && y_pointer == 89)
||(x_pointer == 110 && y_pointer == 89)
||(x_pointer == 111 && y_pointer == 89)
||(x_pointer == 112 && y_pointer == 89)
||(x_pointer == 122 && y_pointer == 89)
||(x_pointer == 123 && y_pointer == 89)
||(x_pointer == 124 && y_pointer == 89)
||(x_pointer == 125 && y_pointer == 89)
||(x_pointer == 126 && y_pointer == 89)
||(x_pointer == 127 && y_pointer == 89)
||(x_pointer == 128 && y_pointer == 89)
||(x_pointer == 129 && y_pointer == 89)
||(x_pointer == 130 && y_pointer == 89)
||(x_pointer == 140 && y_pointer == 89)
||(x_pointer == 141 && y_pointer == 89)
||(x_pointer == 142 && y_pointer == 89)
||(x_pointer == 143 && y_pointer == 89)
||(x_pointer == 144 && y_pointer == 89)
||(x_pointer == 145 && y_pointer == 89)
||(x_pointer == 146 && y_pointer == 89)
||(x_pointer == 147 && y_pointer == 89)
||(x_pointer == 148 && y_pointer == 89)
||(x_pointer == 155 && y_pointer == 89)
||(x_pointer == 156 && y_pointer == 89)
||(x_pointer == 157 && y_pointer == 89)
||(x_pointer == 2 && y_pointer == 90)
||(x_pointer == 3 && y_pointer == 90)
||(x_pointer == 4 && y_pointer == 90)
||(x_pointer == 14 && y_pointer == 90)
||(x_pointer == 15 && y_pointer == 90)
||(x_pointer == 16 && y_pointer == 90)
||(x_pointer == 17 && y_pointer == 90)
||(x_pointer == 18 && y_pointer == 90)
||(x_pointer == 19 && y_pointer == 90)
||(x_pointer == 20 && y_pointer == 90)
||(x_pointer == 21 && y_pointer == 90)
||(x_pointer == 22 && y_pointer == 90)
||(x_pointer == 32 && y_pointer == 90)
||(x_pointer == 33 && y_pointer == 90)
||(x_pointer == 34 && y_pointer == 90)
||(x_pointer == 35 && y_pointer == 90)
||(x_pointer == 36 && y_pointer == 90)
||(x_pointer == 37 && y_pointer == 90)
||(x_pointer == 38 && y_pointer == 90)
||(x_pointer == 39 && y_pointer == 90)
||(x_pointer == 40 && y_pointer == 90)
||(x_pointer == 50 && y_pointer == 90)
||(x_pointer == 51 && y_pointer == 90)
||(x_pointer == 52 && y_pointer == 90)
||(x_pointer == 53 && y_pointer == 90)
||(x_pointer == 54 && y_pointer == 90)
||(x_pointer == 55 && y_pointer == 90)
||(x_pointer == 56 && y_pointer == 90)
||(x_pointer == 57 && y_pointer == 90)
||(x_pointer == 58 && y_pointer == 90)
||(x_pointer == 68 && y_pointer == 90)
||(x_pointer == 69 && y_pointer == 90)
||(x_pointer == 70 && y_pointer == 90)
||(x_pointer == 71 && y_pointer == 90)
||(x_pointer == 72 && y_pointer == 90)
||(x_pointer == 73 && y_pointer == 90)
||(x_pointer == 74 && y_pointer == 90)
||(x_pointer == 75 && y_pointer == 90)
||(x_pointer == 76 && y_pointer == 90)
||(x_pointer == 86 && y_pointer == 90)
||(x_pointer == 87 && y_pointer == 90)
||(x_pointer == 88 && y_pointer == 90)
||(x_pointer == 89 && y_pointer == 90)
||(x_pointer == 90 && y_pointer == 90)
||(x_pointer == 91 && y_pointer == 90)
||(x_pointer == 92 && y_pointer == 90)
||(x_pointer == 93 && y_pointer == 90)
||(x_pointer == 94 && y_pointer == 90)
||(x_pointer == 104 && y_pointer == 90)
||(x_pointer == 105 && y_pointer == 90)
||(x_pointer == 106 && y_pointer == 90)
||(x_pointer == 107 && y_pointer == 90)
||(x_pointer == 108 && y_pointer == 90)
||(x_pointer == 109 && y_pointer == 90)
||(x_pointer == 110 && y_pointer == 90)
||(x_pointer == 111 && y_pointer == 90)
||(x_pointer == 112 && y_pointer == 90)
||(x_pointer == 122 && y_pointer == 90)
||(x_pointer == 123 && y_pointer == 90)
||(x_pointer == 124 && y_pointer == 90)
||(x_pointer == 125 && y_pointer == 90)
||(x_pointer == 126 && y_pointer == 90)
||(x_pointer == 127 && y_pointer == 90)
||(x_pointer == 128 && y_pointer == 90)
||(x_pointer == 129 && y_pointer == 90)
||(x_pointer == 130 && y_pointer == 90)
||(x_pointer == 140 && y_pointer == 90)
||(x_pointer == 141 && y_pointer == 90)
||(x_pointer == 142 && y_pointer == 90)
||(x_pointer == 143 && y_pointer == 90)
||(x_pointer == 144 && y_pointer == 90)
||(x_pointer == 145 && y_pointer == 90)
||(x_pointer == 146 && y_pointer == 90)
||(x_pointer == 147 && y_pointer == 90)
||(x_pointer == 148 && y_pointer == 90)
||(x_pointer == 155 && y_pointer == 90)
||(x_pointer == 156 && y_pointer == 90)
||(x_pointer == 157 && y_pointer == 90)
||(x_pointer == 2 && y_pointer == 91)
||(x_pointer == 3 && y_pointer == 91)
||(x_pointer == 4 && y_pointer == 91)
||(x_pointer == 14 && y_pointer == 91)
||(x_pointer == 15 && y_pointer == 91)
||(x_pointer == 16 && y_pointer == 91)
||(x_pointer == 17 && y_pointer == 91)
||(x_pointer == 18 && y_pointer == 91)
||(x_pointer == 19 && y_pointer == 91)
||(x_pointer == 20 && y_pointer == 91)
||(x_pointer == 21 && y_pointer == 91)
||(x_pointer == 22 && y_pointer == 91)
||(x_pointer == 32 && y_pointer == 91)
||(x_pointer == 33 && y_pointer == 91)
||(x_pointer == 34 && y_pointer == 91)
||(x_pointer == 35 && y_pointer == 91)
||(x_pointer == 36 && y_pointer == 91)
||(x_pointer == 37 && y_pointer == 91)
||(x_pointer == 38 && y_pointer == 91)
||(x_pointer == 39 && y_pointer == 91)
||(x_pointer == 40 && y_pointer == 91)
||(x_pointer == 50 && y_pointer == 91)
||(x_pointer == 51 && y_pointer == 91)
||(x_pointer == 52 && y_pointer == 91)
||(x_pointer == 53 && y_pointer == 91)
||(x_pointer == 54 && y_pointer == 91)
||(x_pointer == 55 && y_pointer == 91)
||(x_pointer == 56 && y_pointer == 91)
||(x_pointer == 57 && y_pointer == 91)
||(x_pointer == 58 && y_pointer == 91)
||(x_pointer == 68 && y_pointer == 91)
||(x_pointer == 69 && y_pointer == 91)
||(x_pointer == 70 && y_pointer == 91)
||(x_pointer == 71 && y_pointer == 91)
||(x_pointer == 72 && y_pointer == 91)
||(x_pointer == 73 && y_pointer == 91)
||(x_pointer == 74 && y_pointer == 91)
||(x_pointer == 75 && y_pointer == 91)
||(x_pointer == 76 && y_pointer == 91)
||(x_pointer == 86 && y_pointer == 91)
||(x_pointer == 87 && y_pointer == 91)
||(x_pointer == 88 && y_pointer == 91)
||(x_pointer == 89 && y_pointer == 91)
||(x_pointer == 90 && y_pointer == 91)
||(x_pointer == 91 && y_pointer == 91)
||(x_pointer == 92 && y_pointer == 91)
||(x_pointer == 93 && y_pointer == 91)
||(x_pointer == 94 && y_pointer == 91)
||(x_pointer == 104 && y_pointer == 91)
||(x_pointer == 105 && y_pointer == 91)
||(x_pointer == 106 && y_pointer == 91)
||(x_pointer == 107 && y_pointer == 91)
||(x_pointer == 108 && y_pointer == 91)
||(x_pointer == 109 && y_pointer == 91)
||(x_pointer == 110 && y_pointer == 91)
||(x_pointer == 111 && y_pointer == 91)
||(x_pointer == 112 && y_pointer == 91)
||(x_pointer == 122 && y_pointer == 91)
||(x_pointer == 123 && y_pointer == 91)
||(x_pointer == 124 && y_pointer == 91)
||(x_pointer == 125 && y_pointer == 91)
||(x_pointer == 126 && y_pointer == 91)
||(x_pointer == 127 && y_pointer == 91)
||(x_pointer == 128 && y_pointer == 91)
||(x_pointer == 129 && y_pointer == 91)
||(x_pointer == 130 && y_pointer == 91)
||(x_pointer == 140 && y_pointer == 91)
||(x_pointer == 141 && y_pointer == 91)
||(x_pointer == 142 && y_pointer == 91)
||(x_pointer == 143 && y_pointer == 91)
||(x_pointer == 144 && y_pointer == 91)
||(x_pointer == 145 && y_pointer == 91)
||(x_pointer == 146 && y_pointer == 91)
||(x_pointer == 147 && y_pointer == 91)
||(x_pointer == 148 && y_pointer == 91)
||(x_pointer == 155 && y_pointer == 91)
||(x_pointer == 156 && y_pointer == 91)
||(x_pointer == 157 && y_pointer == 91)
||(x_pointer == 2 && y_pointer == 92)
||(x_pointer == 3 && y_pointer == 92)
||(x_pointer == 4 && y_pointer == 92)
||(x_pointer == 14 && y_pointer == 92)
||(x_pointer == 15 && y_pointer == 92)
||(x_pointer == 16 && y_pointer == 92)
||(x_pointer == 17 && y_pointer == 92)
||(x_pointer == 18 && y_pointer == 92)
||(x_pointer == 19 && y_pointer == 92)
||(x_pointer == 20 && y_pointer == 92)
||(x_pointer == 21 && y_pointer == 92)
||(x_pointer == 22 && y_pointer == 92)
||(x_pointer == 32 && y_pointer == 92)
||(x_pointer == 33 && y_pointer == 92)
||(x_pointer == 34 && y_pointer == 92)
||(x_pointer == 35 && y_pointer == 92)
||(x_pointer == 36 && y_pointer == 92)
||(x_pointer == 37 && y_pointer == 92)
||(x_pointer == 38 && y_pointer == 92)
||(x_pointer == 39 && y_pointer == 92)
||(x_pointer == 40 && y_pointer == 92)
||(x_pointer == 50 && y_pointer == 92)
||(x_pointer == 51 && y_pointer == 92)
||(x_pointer == 52 && y_pointer == 92)
||(x_pointer == 53 && y_pointer == 92)
||(x_pointer == 54 && y_pointer == 92)
||(x_pointer == 55 && y_pointer == 92)
||(x_pointer == 56 && y_pointer == 92)
||(x_pointer == 57 && y_pointer == 92)
||(x_pointer == 58 && y_pointer == 92)
||(x_pointer == 68 && y_pointer == 92)
||(x_pointer == 69 && y_pointer == 92)
||(x_pointer == 70 && y_pointer == 92)
||(x_pointer == 71 && y_pointer == 92)
||(x_pointer == 72 && y_pointer == 92)
||(x_pointer == 73 && y_pointer == 92)
||(x_pointer == 74 && y_pointer == 92)
||(x_pointer == 75 && y_pointer == 92)
||(x_pointer == 76 && y_pointer == 92)
||(x_pointer == 86 && y_pointer == 92)
||(x_pointer == 87 && y_pointer == 92)
||(x_pointer == 88 && y_pointer == 92)
||(x_pointer == 89 && y_pointer == 92)
||(x_pointer == 90 && y_pointer == 92)
||(x_pointer == 91 && y_pointer == 92)
||(x_pointer == 92 && y_pointer == 92)
||(x_pointer == 93 && y_pointer == 92)
||(x_pointer == 94 && y_pointer == 92)
||(x_pointer == 104 && y_pointer == 92)
||(x_pointer == 105 && y_pointer == 92)
||(x_pointer == 106 && y_pointer == 92)
||(x_pointer == 107 && y_pointer == 92)
||(x_pointer == 108 && y_pointer == 92)
||(x_pointer == 109 && y_pointer == 92)
||(x_pointer == 110 && y_pointer == 92)
||(x_pointer == 111 && y_pointer == 92)
||(x_pointer == 112 && y_pointer == 92)
||(x_pointer == 122 && y_pointer == 92)
||(x_pointer == 123 && y_pointer == 92)
||(x_pointer == 124 && y_pointer == 92)
||(x_pointer == 125 && y_pointer == 92)
||(x_pointer == 126 && y_pointer == 92)
||(x_pointer == 127 && y_pointer == 92)
||(x_pointer == 128 && y_pointer == 92)
||(x_pointer == 129 && y_pointer == 92)
||(x_pointer == 130 && y_pointer == 92)
||(x_pointer == 140 && y_pointer == 92)
||(x_pointer == 141 && y_pointer == 92)
||(x_pointer == 142 && y_pointer == 92)
||(x_pointer == 143 && y_pointer == 92)
||(x_pointer == 144 && y_pointer == 92)
||(x_pointer == 145 && y_pointer == 92)
||(x_pointer == 146 && y_pointer == 92)
||(x_pointer == 147 && y_pointer == 92)
||(x_pointer == 148 && y_pointer == 92)
||(x_pointer == 155 && y_pointer == 92)
||(x_pointer == 156 && y_pointer == 92)
||(x_pointer == 157 && y_pointer == 92)
||(x_pointer == 2 && y_pointer == 93)
||(x_pointer == 3 && y_pointer == 93)
||(x_pointer == 4 && y_pointer == 93)
||(x_pointer == 14 && y_pointer == 93)
||(x_pointer == 15 && y_pointer == 93)
||(x_pointer == 16 && y_pointer == 93)
||(x_pointer == 17 && y_pointer == 93)
||(x_pointer == 18 && y_pointer == 93)
||(x_pointer == 19 && y_pointer == 93)
||(x_pointer == 20 && y_pointer == 93)
||(x_pointer == 21 && y_pointer == 93)
||(x_pointer == 22 && y_pointer == 93)
||(x_pointer == 32 && y_pointer == 93)
||(x_pointer == 33 && y_pointer == 93)
||(x_pointer == 34 && y_pointer == 93)
||(x_pointer == 35 && y_pointer == 93)
||(x_pointer == 36 && y_pointer == 93)
||(x_pointer == 37 && y_pointer == 93)
||(x_pointer == 38 && y_pointer == 93)
||(x_pointer == 39 && y_pointer == 93)
||(x_pointer == 40 && y_pointer == 93)
||(x_pointer == 50 && y_pointer == 93)
||(x_pointer == 51 && y_pointer == 93)
||(x_pointer == 52 && y_pointer == 93)
||(x_pointer == 53 && y_pointer == 93)
||(x_pointer == 54 && y_pointer == 93)
||(x_pointer == 55 && y_pointer == 93)
||(x_pointer == 56 && y_pointer == 93)
||(x_pointer == 57 && y_pointer == 93)
||(x_pointer == 58 && y_pointer == 93)
||(x_pointer == 68 && y_pointer == 93)
||(x_pointer == 69 && y_pointer == 93)
||(x_pointer == 70 && y_pointer == 93)
||(x_pointer == 71 && y_pointer == 93)
||(x_pointer == 72 && y_pointer == 93)
||(x_pointer == 73 && y_pointer == 93)
||(x_pointer == 74 && y_pointer == 93)
||(x_pointer == 75 && y_pointer == 93)
||(x_pointer == 76 && y_pointer == 93)
||(x_pointer == 86 && y_pointer == 93)
||(x_pointer == 87 && y_pointer == 93)
||(x_pointer == 88 && y_pointer == 93)
||(x_pointer == 89 && y_pointer == 93)
||(x_pointer == 90 && y_pointer == 93)
||(x_pointer == 91 && y_pointer == 93)
||(x_pointer == 92 && y_pointer == 93)
||(x_pointer == 93 && y_pointer == 93)
||(x_pointer == 94 && y_pointer == 93)
||(x_pointer == 104 && y_pointer == 93)
||(x_pointer == 105 && y_pointer == 93)
||(x_pointer == 106 && y_pointer == 93)
||(x_pointer == 107 && y_pointer == 93)
||(x_pointer == 108 && y_pointer == 93)
||(x_pointer == 109 && y_pointer == 93)
||(x_pointer == 110 && y_pointer == 93)
||(x_pointer == 111 && y_pointer == 93)
||(x_pointer == 112 && y_pointer == 93)
||(x_pointer == 122 && y_pointer == 93)
||(x_pointer == 123 && y_pointer == 93)
||(x_pointer == 124 && y_pointer == 93)
||(x_pointer == 125 && y_pointer == 93)
||(x_pointer == 126 && y_pointer == 93)
||(x_pointer == 127 && y_pointer == 93)
||(x_pointer == 128 && y_pointer == 93)
||(x_pointer == 129 && y_pointer == 93)
||(x_pointer == 130 && y_pointer == 93)
||(x_pointer == 140 && y_pointer == 93)
||(x_pointer == 141 && y_pointer == 93)
||(x_pointer == 142 && y_pointer == 93)
||(x_pointer == 143 && y_pointer == 93)
||(x_pointer == 144 && y_pointer == 93)
||(x_pointer == 145 && y_pointer == 93)
||(x_pointer == 146 && y_pointer == 93)
||(x_pointer == 147 && y_pointer == 93)
||(x_pointer == 148 && y_pointer == 93)
||(x_pointer == 155 && y_pointer == 93)
||(x_pointer == 156 && y_pointer == 93)
||(x_pointer == 157 && y_pointer == 93)
||(x_pointer == 2 && y_pointer == 94)
||(x_pointer == 3 && y_pointer == 94)
||(x_pointer == 4 && y_pointer == 94)
||(x_pointer == 14 && y_pointer == 94)
||(x_pointer == 15 && y_pointer == 94)
||(x_pointer == 16 && y_pointer == 94)
||(x_pointer == 17 && y_pointer == 94)
||(x_pointer == 18 && y_pointer == 94)
||(x_pointer == 19 && y_pointer == 94)
||(x_pointer == 20 && y_pointer == 94)
||(x_pointer == 21 && y_pointer == 94)
||(x_pointer == 22 && y_pointer == 94)
||(x_pointer == 32 && y_pointer == 94)
||(x_pointer == 33 && y_pointer == 94)
||(x_pointer == 34 && y_pointer == 94)
||(x_pointer == 35 && y_pointer == 94)
||(x_pointer == 36 && y_pointer == 94)
||(x_pointer == 37 && y_pointer == 94)
||(x_pointer == 38 && y_pointer == 94)
||(x_pointer == 39 && y_pointer == 94)
||(x_pointer == 40 && y_pointer == 94)
||(x_pointer == 50 && y_pointer == 94)
||(x_pointer == 51 && y_pointer == 94)
||(x_pointer == 52 && y_pointer == 94)
||(x_pointer == 53 && y_pointer == 94)
||(x_pointer == 54 && y_pointer == 94)
||(x_pointer == 55 && y_pointer == 94)
||(x_pointer == 56 && y_pointer == 94)
||(x_pointer == 57 && y_pointer == 94)
||(x_pointer == 58 && y_pointer == 94)
||(x_pointer == 68 && y_pointer == 94)
||(x_pointer == 69 && y_pointer == 94)
||(x_pointer == 70 && y_pointer == 94)
||(x_pointer == 71 && y_pointer == 94)
||(x_pointer == 72 && y_pointer == 94)
||(x_pointer == 73 && y_pointer == 94)
||(x_pointer == 74 && y_pointer == 94)
||(x_pointer == 75 && y_pointer == 94)
||(x_pointer == 76 && y_pointer == 94)
||(x_pointer == 86 && y_pointer == 94)
||(x_pointer == 87 && y_pointer == 94)
||(x_pointer == 88 && y_pointer == 94)
||(x_pointer == 89 && y_pointer == 94)
||(x_pointer == 90 && y_pointer == 94)
||(x_pointer == 91 && y_pointer == 94)
||(x_pointer == 92 && y_pointer == 94)
||(x_pointer == 93 && y_pointer == 94)
||(x_pointer == 94 && y_pointer == 94)
||(x_pointer == 104 && y_pointer == 94)
||(x_pointer == 105 && y_pointer == 94)
||(x_pointer == 106 && y_pointer == 94)
||(x_pointer == 107 && y_pointer == 94)
||(x_pointer == 108 && y_pointer == 94)
||(x_pointer == 109 && y_pointer == 94)
||(x_pointer == 110 && y_pointer == 94)
||(x_pointer == 111 && y_pointer == 94)
||(x_pointer == 112 && y_pointer == 94)
||(x_pointer == 122 && y_pointer == 94)
||(x_pointer == 123 && y_pointer == 94)
||(x_pointer == 124 && y_pointer == 94)
||(x_pointer == 125 && y_pointer == 94)
||(x_pointer == 126 && y_pointer == 94)
||(x_pointer == 127 && y_pointer == 94)
||(x_pointer == 128 && y_pointer == 94)
||(x_pointer == 129 && y_pointer == 94)
||(x_pointer == 130 && y_pointer == 94)
||(x_pointer == 140 && y_pointer == 94)
||(x_pointer == 141 && y_pointer == 94)
||(x_pointer == 142 && y_pointer == 94)
||(x_pointer == 143 && y_pointer == 94)
||(x_pointer == 144 && y_pointer == 94)
||(x_pointer == 145 && y_pointer == 94)
||(x_pointer == 146 && y_pointer == 94)
||(x_pointer == 147 && y_pointer == 94)
||(x_pointer == 148 && y_pointer == 94)
||(x_pointer == 155 && y_pointer == 94)
||(x_pointer == 156 && y_pointer == 94)
||(x_pointer == 157 && y_pointer == 94)
||(x_pointer == 2 && y_pointer == 95)
||(x_pointer == 3 && y_pointer == 95)
||(x_pointer == 4 && y_pointer == 95)
||(x_pointer == 155 && y_pointer == 95)
||(x_pointer == 156 && y_pointer == 95)
||(x_pointer == 157 && y_pointer == 95)
||(x_pointer == 2 && y_pointer == 96)
||(x_pointer == 3 && y_pointer == 96)
||(x_pointer == 4 && y_pointer == 96)
||(x_pointer == 155 && y_pointer == 96)
||(x_pointer == 156 && y_pointer == 96)
||(x_pointer == 157 && y_pointer == 96)
||(x_pointer == 2 && y_pointer == 97)
||(x_pointer == 3 && y_pointer == 97)
||(x_pointer == 4 && y_pointer == 97)
||(x_pointer == 155 && y_pointer == 97)
||(x_pointer == 156 && y_pointer == 97)
||(x_pointer == 157 && y_pointer == 97)
||(x_pointer == 2 && y_pointer == 98)
||(x_pointer == 3 && y_pointer == 98)
||(x_pointer == 4 && y_pointer == 98)
||(x_pointer == 155 && y_pointer == 98)
||(x_pointer == 156 && y_pointer == 98)
||(x_pointer == 157 && y_pointer == 98)
||(x_pointer == 2 && y_pointer == 99)
||(x_pointer == 3 && y_pointer == 99)
||(x_pointer == 4 && y_pointer == 99)
||(x_pointer == 155 && y_pointer == 99)
||(x_pointer == 156 && y_pointer == 99)
||(x_pointer == 157 && y_pointer == 99)
||(x_pointer == 2 && y_pointer == 100)
||(x_pointer == 3 && y_pointer == 100)
||(x_pointer == 4 && y_pointer == 100)
||(x_pointer == 155 && y_pointer == 100)
||(x_pointer == 156 && y_pointer == 100)
||(x_pointer == 157 && y_pointer == 100)
||(x_pointer == 2 && y_pointer == 101)
||(x_pointer == 3 && y_pointer == 101)
||(x_pointer == 4 && y_pointer == 101)
||(x_pointer == 155 && y_pointer == 101)
||(x_pointer == 156 && y_pointer == 101)
||(x_pointer == 157 && y_pointer == 101)
||(x_pointer == 2 && y_pointer == 102)
||(x_pointer == 3 && y_pointer == 102)
||(x_pointer == 4 && y_pointer == 102)
||(x_pointer == 155 && y_pointer == 102)
||(x_pointer == 156 && y_pointer == 102)
||(x_pointer == 157 && y_pointer == 102)
||(x_pointer == 2 && y_pointer == 103)
||(x_pointer == 3 && y_pointer == 103)
||(x_pointer == 4 && y_pointer == 103)
||(x_pointer == 155 && y_pointer == 103)
||(x_pointer == 156 && y_pointer == 103)
||(x_pointer == 157 && y_pointer == 103)
||(x_pointer == 2 && y_pointer == 104)
||(x_pointer == 3 && y_pointer == 104)
||(x_pointer == 4 && y_pointer == 104)
||(x_pointer == 14 && y_pointer == 104)
||(x_pointer == 15 && y_pointer == 104)
||(x_pointer == 16 && y_pointer == 104)
||(x_pointer == 17 && y_pointer == 104)
||(x_pointer == 18 && y_pointer == 104)
||(x_pointer == 19 && y_pointer == 104)
||(x_pointer == 20 && y_pointer == 104)
||(x_pointer == 21 && y_pointer == 104)
||(x_pointer == 22 && y_pointer == 104)
||(x_pointer == 32 && y_pointer == 104)
||(x_pointer == 33 && y_pointer == 104)
||(x_pointer == 34 && y_pointer == 104)
||(x_pointer == 35 && y_pointer == 104)
||(x_pointer == 36 && y_pointer == 104)
||(x_pointer == 37 && y_pointer == 104)
||(x_pointer == 38 && y_pointer == 104)
||(x_pointer == 39 && y_pointer == 104)
||(x_pointer == 40 && y_pointer == 104)
||(x_pointer == 50 && y_pointer == 104)
||(x_pointer == 51 && y_pointer == 104)
||(x_pointer == 52 && y_pointer == 104)
||(x_pointer == 53 && y_pointer == 104)
||(x_pointer == 54 && y_pointer == 104)
||(x_pointer == 55 && y_pointer == 104)
||(x_pointer == 56 && y_pointer == 104)
||(x_pointer == 57 && y_pointer == 104)
||(x_pointer == 58 && y_pointer == 104)
||(x_pointer == 68 && y_pointer == 104)
||(x_pointer == 69 && y_pointer == 104)
||(x_pointer == 70 && y_pointer == 104)
||(x_pointer == 71 && y_pointer == 104)
||(x_pointer == 72 && y_pointer == 104)
||(x_pointer == 73 && y_pointer == 104)
||(x_pointer == 74 && y_pointer == 104)
||(x_pointer == 75 && y_pointer == 104)
||(x_pointer == 76 && y_pointer == 104)
||(x_pointer == 86 && y_pointer == 104)
||(x_pointer == 87 && y_pointer == 104)
||(x_pointer == 88 && y_pointer == 104)
||(x_pointer == 89 && y_pointer == 104)
||(x_pointer == 90 && y_pointer == 104)
||(x_pointer == 91 && y_pointer == 104)
||(x_pointer == 92 && y_pointer == 104)
||(x_pointer == 93 && y_pointer == 104)
||(x_pointer == 94 && y_pointer == 104)
||(x_pointer == 104 && y_pointer == 104)
||(x_pointer == 105 && y_pointer == 104)
||(x_pointer == 106 && y_pointer == 104)
||(x_pointer == 107 && y_pointer == 104)
||(x_pointer == 108 && y_pointer == 104)
||(x_pointer == 109 && y_pointer == 104)
||(x_pointer == 110 && y_pointer == 104)
||(x_pointer == 111 && y_pointer == 104)
||(x_pointer == 112 && y_pointer == 104)
||(x_pointer == 122 && y_pointer == 104)
||(x_pointer == 123 && y_pointer == 104)
||(x_pointer == 124 && y_pointer == 104)
||(x_pointer == 125 && y_pointer == 104)
||(x_pointer == 126 && y_pointer == 104)
||(x_pointer == 127 && y_pointer == 104)
||(x_pointer == 128 && y_pointer == 104)
||(x_pointer == 129 && y_pointer == 104)
||(x_pointer == 130 && y_pointer == 104)
||(x_pointer == 140 && y_pointer == 104)
||(x_pointer == 141 && y_pointer == 104)
||(x_pointer == 142 && y_pointer == 104)
||(x_pointer == 143 && y_pointer == 104)
||(x_pointer == 144 && y_pointer == 104)
||(x_pointer == 145 && y_pointer == 104)
||(x_pointer == 146 && y_pointer == 104)
||(x_pointer == 147 && y_pointer == 104)
||(x_pointer == 148 && y_pointer == 104)
||(x_pointer == 155 && y_pointer == 104)
||(x_pointer == 156 && y_pointer == 104)
||(x_pointer == 157 && y_pointer == 104)
||(x_pointer == 2 && y_pointer == 105)
||(x_pointer == 3 && y_pointer == 105)
||(x_pointer == 4 && y_pointer == 105)
||(x_pointer == 14 && y_pointer == 105)
||(x_pointer == 15 && y_pointer == 105)
||(x_pointer == 16 && y_pointer == 105)
||(x_pointer == 17 && y_pointer == 105)
||(x_pointer == 18 && y_pointer == 105)
||(x_pointer == 19 && y_pointer == 105)
||(x_pointer == 20 && y_pointer == 105)
||(x_pointer == 21 && y_pointer == 105)
||(x_pointer == 22 && y_pointer == 105)
||(x_pointer == 32 && y_pointer == 105)
||(x_pointer == 33 && y_pointer == 105)
||(x_pointer == 34 && y_pointer == 105)
||(x_pointer == 35 && y_pointer == 105)
||(x_pointer == 36 && y_pointer == 105)
||(x_pointer == 37 && y_pointer == 105)
||(x_pointer == 38 && y_pointer == 105)
||(x_pointer == 39 && y_pointer == 105)
||(x_pointer == 40 && y_pointer == 105)
||(x_pointer == 50 && y_pointer == 105)
||(x_pointer == 51 && y_pointer == 105)
||(x_pointer == 52 && y_pointer == 105)
||(x_pointer == 53 && y_pointer == 105)
||(x_pointer == 54 && y_pointer == 105)
||(x_pointer == 55 && y_pointer == 105)
||(x_pointer == 56 && y_pointer == 105)
||(x_pointer == 57 && y_pointer == 105)
||(x_pointer == 58 && y_pointer == 105)
||(x_pointer == 68 && y_pointer == 105)
||(x_pointer == 69 && y_pointer == 105)
||(x_pointer == 70 && y_pointer == 105)
||(x_pointer == 71 && y_pointer == 105)
||(x_pointer == 72 && y_pointer == 105)
||(x_pointer == 73 && y_pointer == 105)
||(x_pointer == 74 && y_pointer == 105)
||(x_pointer == 75 && y_pointer == 105)
||(x_pointer == 76 && y_pointer == 105)
||(x_pointer == 86 && y_pointer == 105)
||(x_pointer == 87 && y_pointer == 105)
||(x_pointer == 88 && y_pointer == 105)
||(x_pointer == 89 && y_pointer == 105)
||(x_pointer == 90 && y_pointer == 105)
||(x_pointer == 91 && y_pointer == 105)
||(x_pointer == 92 && y_pointer == 105)
||(x_pointer == 93 && y_pointer == 105)
||(x_pointer == 94 && y_pointer == 105)
||(x_pointer == 104 && y_pointer == 105)
||(x_pointer == 105 && y_pointer == 105)
||(x_pointer == 106 && y_pointer == 105)
||(x_pointer == 107 && y_pointer == 105)
||(x_pointer == 108 && y_pointer == 105)
||(x_pointer == 109 && y_pointer == 105)
||(x_pointer == 110 && y_pointer == 105)
||(x_pointer == 111 && y_pointer == 105)
||(x_pointer == 112 && y_pointer == 105)
||(x_pointer == 122 && y_pointer == 105)
||(x_pointer == 123 && y_pointer == 105)
||(x_pointer == 124 && y_pointer == 105)
||(x_pointer == 125 && y_pointer == 105)
||(x_pointer == 126 && y_pointer == 105)
||(x_pointer == 127 && y_pointer == 105)
||(x_pointer == 128 && y_pointer == 105)
||(x_pointer == 129 && y_pointer == 105)
||(x_pointer == 130 && y_pointer == 105)
||(x_pointer == 140 && y_pointer == 105)
||(x_pointer == 141 && y_pointer == 105)
||(x_pointer == 142 && y_pointer == 105)
||(x_pointer == 143 && y_pointer == 105)
||(x_pointer == 144 && y_pointer == 105)
||(x_pointer == 145 && y_pointer == 105)
||(x_pointer == 146 && y_pointer == 105)
||(x_pointer == 147 && y_pointer == 105)
||(x_pointer == 148 && y_pointer == 105)
||(x_pointer == 155 && y_pointer == 105)
||(x_pointer == 156 && y_pointer == 105)
||(x_pointer == 157 && y_pointer == 105)
||(x_pointer == 2 && y_pointer == 106)
||(x_pointer == 3 && y_pointer == 106)
||(x_pointer == 4 && y_pointer == 106)
||(x_pointer == 14 && y_pointer == 106)
||(x_pointer == 15 && y_pointer == 106)
||(x_pointer == 16 && y_pointer == 106)
||(x_pointer == 17 && y_pointer == 106)
||(x_pointer == 18 && y_pointer == 106)
||(x_pointer == 19 && y_pointer == 106)
||(x_pointer == 20 && y_pointer == 106)
||(x_pointer == 21 && y_pointer == 106)
||(x_pointer == 22 && y_pointer == 106)
||(x_pointer == 32 && y_pointer == 106)
||(x_pointer == 33 && y_pointer == 106)
||(x_pointer == 34 && y_pointer == 106)
||(x_pointer == 35 && y_pointer == 106)
||(x_pointer == 36 && y_pointer == 106)
||(x_pointer == 37 && y_pointer == 106)
||(x_pointer == 38 && y_pointer == 106)
||(x_pointer == 39 && y_pointer == 106)
||(x_pointer == 40 && y_pointer == 106)
||(x_pointer == 50 && y_pointer == 106)
||(x_pointer == 51 && y_pointer == 106)
||(x_pointer == 52 && y_pointer == 106)
||(x_pointer == 53 && y_pointer == 106)
||(x_pointer == 54 && y_pointer == 106)
||(x_pointer == 55 && y_pointer == 106)
||(x_pointer == 56 && y_pointer == 106)
||(x_pointer == 57 && y_pointer == 106)
||(x_pointer == 58 && y_pointer == 106)
||(x_pointer == 68 && y_pointer == 106)
||(x_pointer == 69 && y_pointer == 106)
||(x_pointer == 70 && y_pointer == 106)
||(x_pointer == 71 && y_pointer == 106)
||(x_pointer == 72 && y_pointer == 106)
||(x_pointer == 73 && y_pointer == 106)
||(x_pointer == 74 && y_pointer == 106)
||(x_pointer == 75 && y_pointer == 106)
||(x_pointer == 76 && y_pointer == 106)
||(x_pointer == 86 && y_pointer == 106)
||(x_pointer == 87 && y_pointer == 106)
||(x_pointer == 88 && y_pointer == 106)
||(x_pointer == 89 && y_pointer == 106)
||(x_pointer == 90 && y_pointer == 106)
||(x_pointer == 91 && y_pointer == 106)
||(x_pointer == 92 && y_pointer == 106)
||(x_pointer == 93 && y_pointer == 106)
||(x_pointer == 94 && y_pointer == 106)
||(x_pointer == 104 && y_pointer == 106)
||(x_pointer == 105 && y_pointer == 106)
||(x_pointer == 106 && y_pointer == 106)
||(x_pointer == 107 && y_pointer == 106)
||(x_pointer == 108 && y_pointer == 106)
||(x_pointer == 109 && y_pointer == 106)
||(x_pointer == 110 && y_pointer == 106)
||(x_pointer == 111 && y_pointer == 106)
||(x_pointer == 112 && y_pointer == 106)
||(x_pointer == 122 && y_pointer == 106)
||(x_pointer == 123 && y_pointer == 106)
||(x_pointer == 124 && y_pointer == 106)
||(x_pointer == 125 && y_pointer == 106)
||(x_pointer == 126 && y_pointer == 106)
||(x_pointer == 127 && y_pointer == 106)
||(x_pointer == 128 && y_pointer == 106)
||(x_pointer == 129 && y_pointer == 106)
||(x_pointer == 130 && y_pointer == 106)
||(x_pointer == 140 && y_pointer == 106)
||(x_pointer == 141 && y_pointer == 106)
||(x_pointer == 142 && y_pointer == 106)
||(x_pointer == 143 && y_pointer == 106)
||(x_pointer == 144 && y_pointer == 106)
||(x_pointer == 145 && y_pointer == 106)
||(x_pointer == 146 && y_pointer == 106)
||(x_pointer == 147 && y_pointer == 106)
||(x_pointer == 148 && y_pointer == 106)
||(x_pointer == 155 && y_pointer == 106)
||(x_pointer == 156 && y_pointer == 106)
||(x_pointer == 157 && y_pointer == 106)
||(x_pointer == 2 && y_pointer == 107)
||(x_pointer == 3 && y_pointer == 107)
||(x_pointer == 4 && y_pointer == 107)
||(x_pointer == 14 && y_pointer == 107)
||(x_pointer == 15 && y_pointer == 107)
||(x_pointer == 16 && y_pointer == 107)
||(x_pointer == 17 && y_pointer == 107)
||(x_pointer == 18 && y_pointer == 107)
||(x_pointer == 19 && y_pointer == 107)
||(x_pointer == 20 && y_pointer == 107)
||(x_pointer == 21 && y_pointer == 107)
||(x_pointer == 22 && y_pointer == 107)
||(x_pointer == 32 && y_pointer == 107)
||(x_pointer == 33 && y_pointer == 107)
||(x_pointer == 34 && y_pointer == 107)
||(x_pointer == 35 && y_pointer == 107)
||(x_pointer == 36 && y_pointer == 107)
||(x_pointer == 37 && y_pointer == 107)
||(x_pointer == 38 && y_pointer == 107)
||(x_pointer == 39 && y_pointer == 107)
||(x_pointer == 40 && y_pointer == 107)
||(x_pointer == 50 && y_pointer == 107)
||(x_pointer == 51 && y_pointer == 107)
||(x_pointer == 52 && y_pointer == 107)
||(x_pointer == 53 && y_pointer == 107)
||(x_pointer == 54 && y_pointer == 107)
||(x_pointer == 55 && y_pointer == 107)
||(x_pointer == 56 && y_pointer == 107)
||(x_pointer == 57 && y_pointer == 107)
||(x_pointer == 58 && y_pointer == 107)
||(x_pointer == 68 && y_pointer == 107)
||(x_pointer == 69 && y_pointer == 107)
||(x_pointer == 70 && y_pointer == 107)
||(x_pointer == 71 && y_pointer == 107)
||(x_pointer == 72 && y_pointer == 107)
||(x_pointer == 73 && y_pointer == 107)
||(x_pointer == 74 && y_pointer == 107)
||(x_pointer == 75 && y_pointer == 107)
||(x_pointer == 76 && y_pointer == 107)
||(x_pointer == 86 && y_pointer == 107)
||(x_pointer == 87 && y_pointer == 107)
||(x_pointer == 88 && y_pointer == 107)
||(x_pointer == 89 && y_pointer == 107)
||(x_pointer == 90 && y_pointer == 107)
||(x_pointer == 91 && y_pointer == 107)
||(x_pointer == 92 && y_pointer == 107)
||(x_pointer == 93 && y_pointer == 107)
||(x_pointer == 94 && y_pointer == 107)
||(x_pointer == 104 && y_pointer == 107)
||(x_pointer == 105 && y_pointer == 107)
||(x_pointer == 106 && y_pointer == 107)
||(x_pointer == 107 && y_pointer == 107)
||(x_pointer == 108 && y_pointer == 107)
||(x_pointer == 109 && y_pointer == 107)
||(x_pointer == 110 && y_pointer == 107)
||(x_pointer == 111 && y_pointer == 107)
||(x_pointer == 112 && y_pointer == 107)
||(x_pointer == 122 && y_pointer == 107)
||(x_pointer == 123 && y_pointer == 107)
||(x_pointer == 124 && y_pointer == 107)
||(x_pointer == 125 && y_pointer == 107)
||(x_pointer == 126 && y_pointer == 107)
||(x_pointer == 127 && y_pointer == 107)
||(x_pointer == 128 && y_pointer == 107)
||(x_pointer == 129 && y_pointer == 107)
||(x_pointer == 130 && y_pointer == 107)
||(x_pointer == 140 && y_pointer == 107)
||(x_pointer == 141 && y_pointer == 107)
||(x_pointer == 142 && y_pointer == 107)
||(x_pointer == 143 && y_pointer == 107)
||(x_pointer == 144 && y_pointer == 107)
||(x_pointer == 145 && y_pointer == 107)
||(x_pointer == 146 && y_pointer == 107)
||(x_pointer == 147 && y_pointer == 107)
||(x_pointer == 148 && y_pointer == 107)
||(x_pointer == 155 && y_pointer == 107)
||(x_pointer == 156 && y_pointer == 107)
||(x_pointer == 157 && y_pointer == 107)
||(x_pointer == 2 && y_pointer == 108)
||(x_pointer == 3 && y_pointer == 108)
||(x_pointer == 4 && y_pointer == 108)
||(x_pointer == 14 && y_pointer == 108)
||(x_pointer == 15 && y_pointer == 108)
||(x_pointer == 16 && y_pointer == 108)
||(x_pointer == 17 && y_pointer == 108)
||(x_pointer == 18 && y_pointer == 108)
||(x_pointer == 19 && y_pointer == 108)
||(x_pointer == 20 && y_pointer == 108)
||(x_pointer == 21 && y_pointer == 108)
||(x_pointer == 22 && y_pointer == 108)
||(x_pointer == 32 && y_pointer == 108)
||(x_pointer == 33 && y_pointer == 108)
||(x_pointer == 34 && y_pointer == 108)
||(x_pointer == 35 && y_pointer == 108)
||(x_pointer == 36 && y_pointer == 108)
||(x_pointer == 37 && y_pointer == 108)
||(x_pointer == 38 && y_pointer == 108)
||(x_pointer == 39 && y_pointer == 108)
||(x_pointer == 40 && y_pointer == 108)
||(x_pointer == 50 && y_pointer == 108)
||(x_pointer == 51 && y_pointer == 108)
||(x_pointer == 52 && y_pointer == 108)
||(x_pointer == 53 && y_pointer == 108)
||(x_pointer == 54 && y_pointer == 108)
||(x_pointer == 55 && y_pointer == 108)
||(x_pointer == 56 && y_pointer == 108)
||(x_pointer == 57 && y_pointer == 108)
||(x_pointer == 58 && y_pointer == 108)
||(x_pointer == 68 && y_pointer == 108)
||(x_pointer == 69 && y_pointer == 108)
||(x_pointer == 70 && y_pointer == 108)
||(x_pointer == 71 && y_pointer == 108)
||(x_pointer == 72 && y_pointer == 108)
||(x_pointer == 73 && y_pointer == 108)
||(x_pointer == 74 && y_pointer == 108)
||(x_pointer == 75 && y_pointer == 108)
||(x_pointer == 76 && y_pointer == 108)
||(x_pointer == 86 && y_pointer == 108)
||(x_pointer == 87 && y_pointer == 108)
||(x_pointer == 88 && y_pointer == 108)
||(x_pointer == 89 && y_pointer == 108)
||(x_pointer == 90 && y_pointer == 108)
||(x_pointer == 91 && y_pointer == 108)
||(x_pointer == 92 && y_pointer == 108)
||(x_pointer == 93 && y_pointer == 108)
||(x_pointer == 94 && y_pointer == 108)
||(x_pointer == 104 && y_pointer == 108)
||(x_pointer == 105 && y_pointer == 108)
||(x_pointer == 106 && y_pointer == 108)
||(x_pointer == 107 && y_pointer == 108)
||(x_pointer == 108 && y_pointer == 108)
||(x_pointer == 109 && y_pointer == 108)
||(x_pointer == 110 && y_pointer == 108)
||(x_pointer == 111 && y_pointer == 108)
||(x_pointer == 112 && y_pointer == 108)
||(x_pointer == 122 && y_pointer == 108)
||(x_pointer == 123 && y_pointer == 108)
||(x_pointer == 124 && y_pointer == 108)
||(x_pointer == 125 && y_pointer == 108)
||(x_pointer == 126 && y_pointer == 108)
||(x_pointer == 127 && y_pointer == 108)
||(x_pointer == 128 && y_pointer == 108)
||(x_pointer == 129 && y_pointer == 108)
||(x_pointer == 130 && y_pointer == 108)
||(x_pointer == 140 && y_pointer == 108)
||(x_pointer == 141 && y_pointer == 108)
||(x_pointer == 142 && y_pointer == 108)
||(x_pointer == 143 && y_pointer == 108)
||(x_pointer == 144 && y_pointer == 108)
||(x_pointer == 145 && y_pointer == 108)
||(x_pointer == 146 && y_pointer == 108)
||(x_pointer == 147 && y_pointer == 108)
||(x_pointer == 148 && y_pointer == 108)
||(x_pointer == 155 && y_pointer == 108)
||(x_pointer == 156 && y_pointer == 108)
||(x_pointer == 157 && y_pointer == 108)
||(x_pointer == 2 && y_pointer == 109)
||(x_pointer == 3 && y_pointer == 109)
||(x_pointer == 4 && y_pointer == 109)
||(x_pointer == 14 && y_pointer == 109)
||(x_pointer == 15 && y_pointer == 109)
||(x_pointer == 16 && y_pointer == 109)
||(x_pointer == 17 && y_pointer == 109)
||(x_pointer == 18 && y_pointer == 109)
||(x_pointer == 19 && y_pointer == 109)
||(x_pointer == 20 && y_pointer == 109)
||(x_pointer == 21 && y_pointer == 109)
||(x_pointer == 22 && y_pointer == 109)
||(x_pointer == 32 && y_pointer == 109)
||(x_pointer == 33 && y_pointer == 109)
||(x_pointer == 34 && y_pointer == 109)
||(x_pointer == 35 && y_pointer == 109)
||(x_pointer == 36 && y_pointer == 109)
||(x_pointer == 37 && y_pointer == 109)
||(x_pointer == 38 && y_pointer == 109)
||(x_pointer == 39 && y_pointer == 109)
||(x_pointer == 40 && y_pointer == 109)
||(x_pointer == 50 && y_pointer == 109)
||(x_pointer == 51 && y_pointer == 109)
||(x_pointer == 52 && y_pointer == 109)
||(x_pointer == 53 && y_pointer == 109)
||(x_pointer == 54 && y_pointer == 109)
||(x_pointer == 55 && y_pointer == 109)
||(x_pointer == 56 && y_pointer == 109)
||(x_pointer == 57 && y_pointer == 109)
||(x_pointer == 58 && y_pointer == 109)
||(x_pointer == 68 && y_pointer == 109)
||(x_pointer == 69 && y_pointer == 109)
||(x_pointer == 70 && y_pointer == 109)
||(x_pointer == 71 && y_pointer == 109)
||(x_pointer == 72 && y_pointer == 109)
||(x_pointer == 73 && y_pointer == 109)
||(x_pointer == 74 && y_pointer == 109)
||(x_pointer == 75 && y_pointer == 109)
||(x_pointer == 76 && y_pointer == 109)
||(x_pointer == 86 && y_pointer == 109)
||(x_pointer == 87 && y_pointer == 109)
||(x_pointer == 88 && y_pointer == 109)
||(x_pointer == 89 && y_pointer == 109)
||(x_pointer == 90 && y_pointer == 109)
||(x_pointer == 91 && y_pointer == 109)
||(x_pointer == 92 && y_pointer == 109)
||(x_pointer == 93 && y_pointer == 109)
||(x_pointer == 94 && y_pointer == 109)
||(x_pointer == 104 && y_pointer == 109)
||(x_pointer == 105 && y_pointer == 109)
||(x_pointer == 106 && y_pointer == 109)
||(x_pointer == 107 && y_pointer == 109)
||(x_pointer == 108 && y_pointer == 109)
||(x_pointer == 109 && y_pointer == 109)
||(x_pointer == 110 && y_pointer == 109)
||(x_pointer == 111 && y_pointer == 109)
||(x_pointer == 112 && y_pointer == 109)
||(x_pointer == 122 && y_pointer == 109)
||(x_pointer == 123 && y_pointer == 109)
||(x_pointer == 124 && y_pointer == 109)
||(x_pointer == 125 && y_pointer == 109)
||(x_pointer == 126 && y_pointer == 109)
||(x_pointer == 127 && y_pointer == 109)
||(x_pointer == 128 && y_pointer == 109)
||(x_pointer == 129 && y_pointer == 109)
||(x_pointer == 130 && y_pointer == 109)
||(x_pointer == 140 && y_pointer == 109)
||(x_pointer == 141 && y_pointer == 109)
||(x_pointer == 142 && y_pointer == 109)
||(x_pointer == 143 && y_pointer == 109)
||(x_pointer == 144 && y_pointer == 109)
||(x_pointer == 145 && y_pointer == 109)
||(x_pointer == 146 && y_pointer == 109)
||(x_pointer == 147 && y_pointer == 109)
||(x_pointer == 148 && y_pointer == 109)
||(x_pointer == 155 && y_pointer == 109)
||(x_pointer == 156 && y_pointer == 109)
||(x_pointer == 157 && y_pointer == 109)
||(x_pointer == 2 && y_pointer == 110)
||(x_pointer == 3 && y_pointer == 110)
||(x_pointer == 4 && y_pointer == 110)
||(x_pointer == 5 && y_pointer == 110)
||(x_pointer == 6 && y_pointer == 110)
||(x_pointer == 7 && y_pointer == 110)
||(x_pointer == 8 && y_pointer == 110)
||(x_pointer == 9 && y_pointer == 110)
||(x_pointer == 10 && y_pointer == 110)
||(x_pointer == 11 && y_pointer == 110)
||(x_pointer == 12 && y_pointer == 110)
||(x_pointer == 13 && y_pointer == 110)
||(x_pointer == 14 && y_pointer == 110)
||(x_pointer == 15 && y_pointer == 110)
||(x_pointer == 16 && y_pointer == 110)
||(x_pointer == 17 && y_pointer == 110)
||(x_pointer == 18 && y_pointer == 110)
||(x_pointer == 19 && y_pointer == 110)
||(x_pointer == 20 && y_pointer == 110)
||(x_pointer == 21 && y_pointer == 110)
||(x_pointer == 22 && y_pointer == 110)
||(x_pointer == 23 && y_pointer == 110)
||(x_pointer == 24 && y_pointer == 110)
||(x_pointer == 25 && y_pointer == 110)
||(x_pointer == 26 && y_pointer == 110)
||(x_pointer == 27 && y_pointer == 110)
||(x_pointer == 28 && y_pointer == 110)
||(x_pointer == 29 && y_pointer == 110)
||(x_pointer == 30 && y_pointer == 110)
||(x_pointer == 31 && y_pointer == 110)
||(x_pointer == 32 && y_pointer == 110)
||(x_pointer == 33 && y_pointer == 110)
||(x_pointer == 34 && y_pointer == 110)
||(x_pointer == 35 && y_pointer == 110)
||(x_pointer == 36 && y_pointer == 110)
||(x_pointer == 37 && y_pointer == 110)
||(x_pointer == 38 && y_pointer == 110)
||(x_pointer == 39 && y_pointer == 110)
||(x_pointer == 40 && y_pointer == 110)
||(x_pointer == 41 && y_pointer == 110)
||(x_pointer == 42 && y_pointer == 110)
||(x_pointer == 43 && y_pointer == 110)
||(x_pointer == 44 && y_pointer == 110)
||(x_pointer == 45 && y_pointer == 110)
||(x_pointer == 46 && y_pointer == 110)
||(x_pointer == 47 && y_pointer == 110)
||(x_pointer == 48 && y_pointer == 110)
||(x_pointer == 49 && y_pointer == 110)
||(x_pointer == 50 && y_pointer == 110)
||(x_pointer == 51 && y_pointer == 110)
||(x_pointer == 52 && y_pointer == 110)
||(x_pointer == 53 && y_pointer == 110)
||(x_pointer == 54 && y_pointer == 110)
||(x_pointer == 55 && y_pointer == 110)
||(x_pointer == 56 && y_pointer == 110)
||(x_pointer == 57 && y_pointer == 110)
||(x_pointer == 58 && y_pointer == 110)
||(x_pointer == 59 && y_pointer == 110)
||(x_pointer == 60 && y_pointer == 110)
||(x_pointer == 61 && y_pointer == 110)
||(x_pointer == 62 && y_pointer == 110)
||(x_pointer == 63 && y_pointer == 110)
||(x_pointer == 64 && y_pointer == 110)
||(x_pointer == 65 && y_pointer == 110)
||(x_pointer == 66 && y_pointer == 110)
||(x_pointer == 67 && y_pointer == 110)
||(x_pointer == 68 && y_pointer == 110)
||(x_pointer == 69 && y_pointer == 110)
||(x_pointer == 70 && y_pointer == 110)
||(x_pointer == 71 && y_pointer == 110)
||(x_pointer == 72 && y_pointer == 110)
||(x_pointer == 73 && y_pointer == 110)
||(x_pointer == 74 && y_pointer == 110)
||(x_pointer == 75 && y_pointer == 110)
||(x_pointer == 76 && y_pointer == 110)
||(x_pointer == 77 && y_pointer == 110)
||(x_pointer == 78 && y_pointer == 110)
||(x_pointer == 79 && y_pointer == 110)
||(x_pointer == 80 && y_pointer == 110)
||(x_pointer == 81 && y_pointer == 110)
||(x_pointer == 82 && y_pointer == 110)
||(x_pointer == 83 && y_pointer == 110)
||(x_pointer == 84 && y_pointer == 110)
||(x_pointer == 85 && y_pointer == 110)
||(x_pointer == 86 && y_pointer == 110)
||(x_pointer == 87 && y_pointer == 110)
||(x_pointer == 88 && y_pointer == 110)
||(x_pointer == 89 && y_pointer == 110)
||(x_pointer == 90 && y_pointer == 110)
||(x_pointer == 91 && y_pointer == 110)
||(x_pointer == 92 && y_pointer == 110)
||(x_pointer == 93 && y_pointer == 110)
||(x_pointer == 94 && y_pointer == 110)
||(x_pointer == 95 && y_pointer == 110)
||(x_pointer == 96 && y_pointer == 110)
||(x_pointer == 97 && y_pointer == 110)
||(x_pointer == 98 && y_pointer == 110)
||(x_pointer == 99 && y_pointer == 110)
||(x_pointer == 100 && y_pointer == 110)
||(x_pointer == 101 && y_pointer == 110)
||(x_pointer == 102 && y_pointer == 110)
||(x_pointer == 103 && y_pointer == 110)
||(x_pointer == 104 && y_pointer == 110)
||(x_pointer == 105 && y_pointer == 110)
||(x_pointer == 106 && y_pointer == 110)
||(x_pointer == 107 && y_pointer == 110)
||(x_pointer == 108 && y_pointer == 110)
||(x_pointer == 109 && y_pointer == 110)
||(x_pointer == 110 && y_pointer == 110)
||(x_pointer == 111 && y_pointer == 110)
||(x_pointer == 112 && y_pointer == 110)
||(x_pointer == 113 && y_pointer == 110)
||(x_pointer == 114 && y_pointer == 110)
||(x_pointer == 115 && y_pointer == 110)
||(x_pointer == 116 && y_pointer == 110)
||(x_pointer == 117 && y_pointer == 110)
||(x_pointer == 118 && y_pointer == 110)
||(x_pointer == 119 && y_pointer == 110)
||(x_pointer == 120 && y_pointer == 110)
||(x_pointer == 121 && y_pointer == 110)
||(x_pointer == 122 && y_pointer == 110)
||(x_pointer == 123 && y_pointer == 110)
||(x_pointer == 124 && y_pointer == 110)
||(x_pointer == 125 && y_pointer == 110)
||(x_pointer == 126 && y_pointer == 110)
||(x_pointer == 127 && y_pointer == 110)
||(x_pointer == 128 && y_pointer == 110)
||(x_pointer == 129 && y_pointer == 110)
||(x_pointer == 130 && y_pointer == 110)
||(x_pointer == 131 && y_pointer == 110)
||(x_pointer == 132 && y_pointer == 110)
||(x_pointer == 133 && y_pointer == 110)
||(x_pointer == 134 && y_pointer == 110)
||(x_pointer == 135 && y_pointer == 110)
||(x_pointer == 136 && y_pointer == 110)
||(x_pointer == 137 && y_pointer == 110)
||(x_pointer == 138 && y_pointer == 110)
||(x_pointer == 139 && y_pointer == 110)
||(x_pointer == 140 && y_pointer == 110)
||(x_pointer == 141 && y_pointer == 110)
||(x_pointer == 142 && y_pointer == 110)
||(x_pointer == 143 && y_pointer == 110)
||(x_pointer == 144 && y_pointer == 110)
||(x_pointer == 145 && y_pointer == 110)
||(x_pointer == 146 && y_pointer == 110)
||(x_pointer == 147 && y_pointer == 110)
||(x_pointer == 148 && y_pointer == 110)
||(x_pointer == 149 && y_pointer == 110)
||(x_pointer == 150 && y_pointer == 110)
||(x_pointer == 151 && y_pointer == 110)
||(x_pointer == 152 && y_pointer == 110)
||(x_pointer == 153 && y_pointer == 110)
||(x_pointer == 154 && y_pointer == 110)
||(x_pointer == 155 && y_pointer == 110)
||(x_pointer == 156 && y_pointer == 110)
||(x_pointer == 157 && y_pointer == 110)
||(x_pointer == 2 && y_pointer == 111)
||(x_pointer == 3 && y_pointer == 111)
||(x_pointer == 4 && y_pointer == 111)
||(x_pointer == 5 && y_pointer == 111)
||(x_pointer == 6 && y_pointer == 111)
||(x_pointer == 7 && y_pointer == 111)
||(x_pointer == 8 && y_pointer == 111)
||(x_pointer == 9 && y_pointer == 111)
||(x_pointer == 10 && y_pointer == 111)
||(x_pointer == 11 && y_pointer == 111)
||(x_pointer == 12 && y_pointer == 111)
||(x_pointer == 13 && y_pointer == 111)
||(x_pointer == 14 && y_pointer == 111)
||(x_pointer == 15 && y_pointer == 111)
||(x_pointer == 16 && y_pointer == 111)
||(x_pointer == 17 && y_pointer == 111)
||(x_pointer == 18 && y_pointer == 111)
||(x_pointer == 19 && y_pointer == 111)
||(x_pointer == 20 && y_pointer == 111)
||(x_pointer == 21 && y_pointer == 111)
||(x_pointer == 22 && y_pointer == 111)
||(x_pointer == 23 && y_pointer == 111)
||(x_pointer == 24 && y_pointer == 111)
||(x_pointer == 25 && y_pointer == 111)
||(x_pointer == 26 && y_pointer == 111)
||(x_pointer == 27 && y_pointer == 111)
||(x_pointer == 28 && y_pointer == 111)
||(x_pointer == 29 && y_pointer == 111)
||(x_pointer == 30 && y_pointer == 111)
||(x_pointer == 31 && y_pointer == 111)
||(x_pointer == 32 && y_pointer == 111)
||(x_pointer == 33 && y_pointer == 111)
||(x_pointer == 34 && y_pointer == 111)
||(x_pointer == 35 && y_pointer == 111)
||(x_pointer == 36 && y_pointer == 111)
||(x_pointer == 37 && y_pointer == 111)
||(x_pointer == 38 && y_pointer == 111)
||(x_pointer == 39 && y_pointer == 111)
||(x_pointer == 40 && y_pointer == 111)
||(x_pointer == 41 && y_pointer == 111)
||(x_pointer == 42 && y_pointer == 111)
||(x_pointer == 43 && y_pointer == 111)
||(x_pointer == 44 && y_pointer == 111)
||(x_pointer == 45 && y_pointer == 111)
||(x_pointer == 46 && y_pointer == 111)
||(x_pointer == 47 && y_pointer == 111)
||(x_pointer == 48 && y_pointer == 111)
||(x_pointer == 49 && y_pointer == 111)
||(x_pointer == 50 && y_pointer == 111)
||(x_pointer == 51 && y_pointer == 111)
||(x_pointer == 52 && y_pointer == 111)
||(x_pointer == 53 && y_pointer == 111)
||(x_pointer == 54 && y_pointer == 111)
||(x_pointer == 55 && y_pointer == 111)
||(x_pointer == 56 && y_pointer == 111)
||(x_pointer == 57 && y_pointer == 111)
||(x_pointer == 58 && y_pointer == 111)
||(x_pointer == 59 && y_pointer == 111)
||(x_pointer == 60 && y_pointer == 111)
||(x_pointer == 61 && y_pointer == 111)
||(x_pointer == 62 && y_pointer == 111)
||(x_pointer == 63 && y_pointer == 111)
||(x_pointer == 64 && y_pointer == 111)
||(x_pointer == 65 && y_pointer == 111)
||(x_pointer == 66 && y_pointer == 111)
||(x_pointer == 67 && y_pointer == 111)
||(x_pointer == 68 && y_pointer == 111)
||(x_pointer == 69 && y_pointer == 111)
||(x_pointer == 70 && y_pointer == 111)
||(x_pointer == 71 && y_pointer == 111)
||(x_pointer == 72 && y_pointer == 111)
||(x_pointer == 73 && y_pointer == 111)
||(x_pointer == 74 && y_pointer == 111)
||(x_pointer == 75 && y_pointer == 111)
||(x_pointer == 76 && y_pointer == 111)
||(x_pointer == 77 && y_pointer == 111)
||(x_pointer == 78 && y_pointer == 111)
||(x_pointer == 79 && y_pointer == 111)
||(x_pointer == 80 && y_pointer == 111)
||(x_pointer == 81 && y_pointer == 111)
||(x_pointer == 82 && y_pointer == 111)
||(x_pointer == 83 && y_pointer == 111)
||(x_pointer == 84 && y_pointer == 111)
||(x_pointer == 85 && y_pointer == 111)
||(x_pointer == 86 && y_pointer == 111)
||(x_pointer == 87 && y_pointer == 111)
||(x_pointer == 88 && y_pointer == 111)
||(x_pointer == 89 && y_pointer == 111)
||(x_pointer == 90 && y_pointer == 111)
||(x_pointer == 91 && y_pointer == 111)
||(x_pointer == 92 && y_pointer == 111)
||(x_pointer == 93 && y_pointer == 111)
||(x_pointer == 94 && y_pointer == 111)
||(x_pointer == 95 && y_pointer == 111)
||(x_pointer == 96 && y_pointer == 111)
||(x_pointer == 97 && y_pointer == 111)
||(x_pointer == 98 && y_pointer == 111)
||(x_pointer == 99 && y_pointer == 111)
||(x_pointer == 100 && y_pointer == 111)
||(x_pointer == 101 && y_pointer == 111)
||(x_pointer == 102 && y_pointer == 111)
||(x_pointer == 103 && y_pointer == 111)
||(x_pointer == 104 && y_pointer == 111)
||(x_pointer == 105 && y_pointer == 111)
||(x_pointer == 106 && y_pointer == 111)
||(x_pointer == 107 && y_pointer == 111)
||(x_pointer == 108 && y_pointer == 111)
||(x_pointer == 109 && y_pointer == 111)
||(x_pointer == 110 && y_pointer == 111)
||(x_pointer == 111 && y_pointer == 111)
||(x_pointer == 112 && y_pointer == 111)
||(x_pointer == 113 && y_pointer == 111)
||(x_pointer == 114 && y_pointer == 111)
||(x_pointer == 115 && y_pointer == 111)
||(x_pointer == 116 && y_pointer == 111)
||(x_pointer == 117 && y_pointer == 111)
||(x_pointer == 118 && y_pointer == 111)
||(x_pointer == 119 && y_pointer == 111)
||(x_pointer == 120 && y_pointer == 111)
||(x_pointer == 121 && y_pointer == 111)
||(x_pointer == 122 && y_pointer == 111)
||(x_pointer == 123 && y_pointer == 111)
||(x_pointer == 124 && y_pointer == 111)
||(x_pointer == 125 && y_pointer == 111)
||(x_pointer == 126 && y_pointer == 111)
||(x_pointer == 127 && y_pointer == 111)
||(x_pointer == 128 && y_pointer == 111)
||(x_pointer == 129 && y_pointer == 111)
||(x_pointer == 130 && y_pointer == 111)
||(x_pointer == 131 && y_pointer == 111)
||(x_pointer == 132 && y_pointer == 111)
||(x_pointer == 133 && y_pointer == 111)
||(x_pointer == 134 && y_pointer == 111)
||(x_pointer == 135 && y_pointer == 111)
||(x_pointer == 136 && y_pointer == 111)
||(x_pointer == 137 && y_pointer == 111)
||(x_pointer == 138 && y_pointer == 111)
||(x_pointer == 139 && y_pointer == 111)
||(x_pointer == 140 && y_pointer == 111)
||(x_pointer == 141 && y_pointer == 111)
||(x_pointer == 142 && y_pointer == 111)
||(x_pointer == 143 && y_pointer == 111)
||(x_pointer == 144 && y_pointer == 111)
||(x_pointer == 145 && y_pointer == 111)
||(x_pointer == 146 && y_pointer == 111)
||(x_pointer == 147 && y_pointer == 111)
||(x_pointer == 148 && y_pointer == 111)
||(x_pointer == 149 && y_pointer == 111)
||(x_pointer == 150 && y_pointer == 111)
||(x_pointer == 151 && y_pointer == 111)
||(x_pointer == 152 && y_pointer == 111)
||(x_pointer == 153 && y_pointer == 111)
||(x_pointer == 154 && y_pointer == 111)
||(x_pointer == 155 && y_pointer == 111)
||(x_pointer == 156 && y_pointer == 111)
||(x_pointer == 157 && y_pointer == 111)
||(x_pointer == 2 && y_pointer == 112)
||(x_pointer == 3 && y_pointer == 112)
||(x_pointer == 4 && y_pointer == 112)
||(x_pointer == 5 && y_pointer == 112)
||(x_pointer == 6 && y_pointer == 112)
||(x_pointer == 7 && y_pointer == 112)
||(x_pointer == 8 && y_pointer == 112)
||(x_pointer == 9 && y_pointer == 112)
||(x_pointer == 10 && y_pointer == 112)
||(x_pointer == 11 && y_pointer == 112)
||(x_pointer == 12 && y_pointer == 112)
||(x_pointer == 13 && y_pointer == 112)
||(x_pointer == 14 && y_pointer == 112)
||(x_pointer == 15 && y_pointer == 112)
||(x_pointer == 16 && y_pointer == 112)
||(x_pointer == 17 && y_pointer == 112)
||(x_pointer == 18 && y_pointer == 112)
||(x_pointer == 19 && y_pointer == 112)
||(x_pointer == 20 && y_pointer == 112)
||(x_pointer == 21 && y_pointer == 112)
||(x_pointer == 22 && y_pointer == 112)
||(x_pointer == 23 && y_pointer == 112)
||(x_pointer == 24 && y_pointer == 112)
||(x_pointer == 25 && y_pointer == 112)
||(x_pointer == 26 && y_pointer == 112)
||(x_pointer == 27 && y_pointer == 112)
||(x_pointer == 28 && y_pointer == 112)
||(x_pointer == 29 && y_pointer == 112)
||(x_pointer == 30 && y_pointer == 112)
||(x_pointer == 31 && y_pointer == 112)
||(x_pointer == 32 && y_pointer == 112)
||(x_pointer == 33 && y_pointer == 112)
||(x_pointer == 34 && y_pointer == 112)
||(x_pointer == 35 && y_pointer == 112)
||(x_pointer == 36 && y_pointer == 112)
||(x_pointer == 37 && y_pointer == 112)
||(x_pointer == 38 && y_pointer == 112)
||(x_pointer == 39 && y_pointer == 112)
||(x_pointer == 40 && y_pointer == 112)
||(x_pointer == 41 && y_pointer == 112)
||(x_pointer == 42 && y_pointer == 112)
||(x_pointer == 43 && y_pointer == 112)
||(x_pointer == 44 && y_pointer == 112)
||(x_pointer == 45 && y_pointer == 112)
||(x_pointer == 46 && y_pointer == 112)
||(x_pointer == 47 && y_pointer == 112)
||(x_pointer == 48 && y_pointer == 112)
||(x_pointer == 49 && y_pointer == 112)
||(x_pointer == 50 && y_pointer == 112)
||(x_pointer == 51 && y_pointer == 112)
||(x_pointer == 52 && y_pointer == 112)
||(x_pointer == 53 && y_pointer == 112)
||(x_pointer == 54 && y_pointer == 112)
||(x_pointer == 55 && y_pointer == 112)
||(x_pointer == 56 && y_pointer == 112)
||(x_pointer == 57 && y_pointer == 112)
||(x_pointer == 58 && y_pointer == 112)
||(x_pointer == 59 && y_pointer == 112)
||(x_pointer == 60 && y_pointer == 112)
||(x_pointer == 61 && y_pointer == 112)
||(x_pointer == 62 && y_pointer == 112)
||(x_pointer == 63 && y_pointer == 112)
||(x_pointer == 64 && y_pointer == 112)
||(x_pointer == 65 && y_pointer == 112)
||(x_pointer == 66 && y_pointer == 112)
||(x_pointer == 67 && y_pointer == 112)
||(x_pointer == 68 && y_pointer == 112)
||(x_pointer == 69 && y_pointer == 112)
||(x_pointer == 70 && y_pointer == 112)
||(x_pointer == 71 && y_pointer == 112)
||(x_pointer == 72 && y_pointer == 112)
||(x_pointer == 73 && y_pointer == 112)
||(x_pointer == 74 && y_pointer == 112)
||(x_pointer == 75 && y_pointer == 112)
||(x_pointer == 76 && y_pointer == 112)
||(x_pointer == 77 && y_pointer == 112)
||(x_pointer == 78 && y_pointer == 112)
||(x_pointer == 79 && y_pointer == 112)
||(x_pointer == 80 && y_pointer == 112)
||(x_pointer == 81 && y_pointer == 112)
||(x_pointer == 82 && y_pointer == 112)
||(x_pointer == 83 && y_pointer == 112)
||(x_pointer == 84 && y_pointer == 112)
||(x_pointer == 85 && y_pointer == 112)
||(x_pointer == 86 && y_pointer == 112)
||(x_pointer == 87 && y_pointer == 112)
||(x_pointer == 88 && y_pointer == 112)
||(x_pointer == 89 && y_pointer == 112)
||(x_pointer == 90 && y_pointer == 112)
||(x_pointer == 91 && y_pointer == 112)
||(x_pointer == 92 && y_pointer == 112)
||(x_pointer == 93 && y_pointer == 112)
||(x_pointer == 94 && y_pointer == 112)
||(x_pointer == 95 && y_pointer == 112)
||(x_pointer == 96 && y_pointer == 112)
||(x_pointer == 97 && y_pointer == 112)
||(x_pointer == 98 && y_pointer == 112)
||(x_pointer == 99 && y_pointer == 112)
||(x_pointer == 100 && y_pointer == 112)
||(x_pointer == 101 && y_pointer == 112)
||(x_pointer == 102 && y_pointer == 112)
||(x_pointer == 103 && y_pointer == 112)
||(x_pointer == 104 && y_pointer == 112)
||(x_pointer == 105 && y_pointer == 112)
||(x_pointer == 106 && y_pointer == 112)
||(x_pointer == 107 && y_pointer == 112)
||(x_pointer == 108 && y_pointer == 112)
||(x_pointer == 109 && y_pointer == 112)
||(x_pointer == 110 && y_pointer == 112)
||(x_pointer == 111 && y_pointer == 112)
||(x_pointer == 112 && y_pointer == 112)
||(x_pointer == 113 && y_pointer == 112)
||(x_pointer == 114 && y_pointer == 112)
||(x_pointer == 115 && y_pointer == 112)
||(x_pointer == 116 && y_pointer == 112)
||(x_pointer == 117 && y_pointer == 112)
||(x_pointer == 118 && y_pointer == 112)
||(x_pointer == 119 && y_pointer == 112)
||(x_pointer == 120 && y_pointer == 112)
||(x_pointer == 121 && y_pointer == 112)
||(x_pointer == 122 && y_pointer == 112)
||(x_pointer == 123 && y_pointer == 112)
||(x_pointer == 124 && y_pointer == 112)
||(x_pointer == 125 && y_pointer == 112)
||(x_pointer == 126 && y_pointer == 112)
||(x_pointer == 127 && y_pointer == 112)
||(x_pointer == 128 && y_pointer == 112)
||(x_pointer == 129 && y_pointer == 112)
||(x_pointer == 130 && y_pointer == 112)
||(x_pointer == 131 && y_pointer == 112)
||(x_pointer == 132 && y_pointer == 112)
||(x_pointer == 133 && y_pointer == 112)
||(x_pointer == 134 && y_pointer == 112)
||(x_pointer == 135 && y_pointer == 112)
||(x_pointer == 136 && y_pointer == 112)
||(x_pointer == 137 && y_pointer == 112)
||(x_pointer == 138 && y_pointer == 112)
||(x_pointer == 139 && y_pointer == 112)
||(x_pointer == 140 && y_pointer == 112)
||(x_pointer == 141 && y_pointer == 112)
||(x_pointer == 142 && y_pointer == 112)
||(x_pointer == 143 && y_pointer == 112)
||(x_pointer == 144 && y_pointer == 112)
||(x_pointer == 145 && y_pointer == 112)
||(x_pointer == 146 && y_pointer == 112)
||(x_pointer == 147 && y_pointer == 112)
||(x_pointer == 148 && y_pointer == 112)
||(x_pointer == 149 && y_pointer == 112)
||(x_pointer == 150 && y_pointer == 112)
||(x_pointer == 151 && y_pointer == 112)
||(x_pointer == 152 && y_pointer == 112)
||(x_pointer == 153 && y_pointer == 112)
||(x_pointer == 154 && y_pointer == 112)
||(x_pointer == 155 && y_pointer == 112)
||(x_pointer == 156 && y_pointer == 112)
||(x_pointer == 157 && y_pointer == 112));
	
	wire barrier_pixel_6 = current_level == 6 && ((x_pointer == 14 && y_pointer == 17)
||(x_pointer == 15 && y_pointer == 17)
||(x_pointer == 16 && y_pointer == 17)
||(x_pointer == 26 && y_pointer == 17)
||(x_pointer == 27 && y_pointer == 17)
||(x_pointer == 28 && y_pointer == 17)
||(x_pointer == 29 && y_pointer == 17)
||(x_pointer == 30 && y_pointer == 17)
||(x_pointer == 31 && y_pointer == 17)
||(x_pointer == 32 && y_pointer == 17)
||(x_pointer == 33 && y_pointer == 17)
||(x_pointer == 34 && y_pointer == 17)
||(x_pointer == 35 && y_pointer == 17)
||(x_pointer == 36 && y_pointer == 17)
||(x_pointer == 37 && y_pointer == 17)
||(x_pointer == 38 && y_pointer == 17)
||(x_pointer == 39 && y_pointer == 17)
||(x_pointer == 40 && y_pointer == 17)
||(x_pointer == 41 && y_pointer == 17)
||(x_pointer == 42 && y_pointer == 17)
||(x_pointer == 43 && y_pointer == 17)
||(x_pointer == 53 && y_pointer == 17)
||(x_pointer == 54 && y_pointer == 17)
||(x_pointer == 55 && y_pointer == 17)
||(x_pointer == 56 && y_pointer == 17)
||(x_pointer == 57 && y_pointer == 17)
||(x_pointer == 58 && y_pointer == 17)
||(x_pointer == 68 && y_pointer == 17)
||(x_pointer == 69 && y_pointer == 17)
||(x_pointer == 70 && y_pointer == 17)
||(x_pointer == 71 && y_pointer == 17)
||(x_pointer == 72 && y_pointer == 17)
||(x_pointer == 73 && y_pointer == 17)
||(x_pointer == 74 && y_pointer == 17)
||(x_pointer == 75 && y_pointer == 17)
||(x_pointer == 76 && y_pointer == 17)
||(x_pointer == 77 && y_pointer == 17)
||(x_pointer == 78 && y_pointer == 17)
||(x_pointer == 79 && y_pointer == 17)
||(x_pointer == 80 && y_pointer == 17)
||(x_pointer == 81 && y_pointer == 17)
||(x_pointer == 82 && y_pointer == 17)
||(x_pointer == 83 && y_pointer == 17)
||(x_pointer == 84 && y_pointer == 17)
||(x_pointer == 85 && y_pointer == 17)
||(x_pointer == 86 && y_pointer == 17)
||(x_pointer == 87 && y_pointer == 17)
||(x_pointer == 88 && y_pointer == 17)
||(x_pointer == 89 && y_pointer == 17)
||(x_pointer == 90 && y_pointer == 17)
||(x_pointer == 91 && y_pointer == 17)
||(x_pointer == 92 && y_pointer == 17)
||(x_pointer == 93 && y_pointer == 17)
||(x_pointer == 94 && y_pointer == 17)
||(x_pointer == 95 && y_pointer == 17)
||(x_pointer == 96 && y_pointer == 17)
||(x_pointer == 97 && y_pointer == 17)
||(x_pointer == 98 && y_pointer == 17)
||(x_pointer == 99 && y_pointer == 17)
||(x_pointer == 100 && y_pointer == 17)
||(x_pointer == 101 && y_pointer == 17)
||(x_pointer == 102 && y_pointer == 17)
||(x_pointer == 103 && y_pointer == 17)
||(x_pointer == 104 && y_pointer == 17)
||(x_pointer == 105 && y_pointer == 17)
||(x_pointer == 106 && y_pointer == 17)
||(x_pointer == 107 && y_pointer == 17)
||(x_pointer == 108 && y_pointer == 17)
||(x_pointer == 109 && y_pointer == 17)
||(x_pointer == 110 && y_pointer == 17)
||(x_pointer == 111 && y_pointer == 17)
||(x_pointer == 112 && y_pointer == 17)
||(x_pointer == 113 && y_pointer == 17)
||(x_pointer == 114 && y_pointer == 17)
||(x_pointer == 115 && y_pointer == 17)
||(x_pointer == 116 && y_pointer == 17)
||(x_pointer == 117 && y_pointer == 17)
||(x_pointer == 118 && y_pointer == 17)
||(x_pointer == 119 && y_pointer == 17)
||(x_pointer == 120 && y_pointer == 17)
||(x_pointer == 121 && y_pointer == 17)
||(x_pointer == 122 && y_pointer == 17)
||(x_pointer == 123 && y_pointer == 17)
||(x_pointer == 124 && y_pointer == 17)
||(x_pointer == 125 && y_pointer == 17)
||(x_pointer == 126 && y_pointer == 17)
||(x_pointer == 127 && y_pointer == 17)
||(x_pointer == 128 && y_pointer == 17)
||(x_pointer == 129 && y_pointer == 17)
||(x_pointer == 130 && y_pointer == 17)
||(x_pointer == 131 && y_pointer == 17)
||(x_pointer == 132 && y_pointer == 17)
||(x_pointer == 133 && y_pointer == 17)
||(x_pointer == 134 && y_pointer == 17)
||(x_pointer == 135 && y_pointer == 17)
||(x_pointer == 136 && y_pointer == 17)
||(x_pointer == 137 && y_pointer == 17)
||(x_pointer == 138 && y_pointer == 17)
||(x_pointer == 139 && y_pointer == 17)
||(x_pointer == 140 && y_pointer == 17)
||(x_pointer == 141 && y_pointer == 17)
||(x_pointer == 142 && y_pointer == 17)
||(x_pointer == 143 && y_pointer == 17)
||(x_pointer == 144 && y_pointer == 17)
||(x_pointer == 145 && y_pointer == 17)
||(x_pointer == 14 && y_pointer == 18)
||(x_pointer == 15 && y_pointer == 18)
||(x_pointer == 16 && y_pointer == 18)
||(x_pointer == 26 && y_pointer == 18)
||(x_pointer == 27 && y_pointer == 18)
||(x_pointer == 28 && y_pointer == 18)
||(x_pointer == 29 && y_pointer == 18)
||(x_pointer == 30 && y_pointer == 18)
||(x_pointer == 31 && y_pointer == 18)
||(x_pointer == 32 && y_pointer == 18)
||(x_pointer == 33 && y_pointer == 18)
||(x_pointer == 34 && y_pointer == 18)
||(x_pointer == 35 && y_pointer == 18)
||(x_pointer == 36 && y_pointer == 18)
||(x_pointer == 37 && y_pointer == 18)
||(x_pointer == 38 && y_pointer == 18)
||(x_pointer == 39 && y_pointer == 18)
||(x_pointer == 40 && y_pointer == 18)
||(x_pointer == 41 && y_pointer == 18)
||(x_pointer == 42 && y_pointer == 18)
||(x_pointer == 43 && y_pointer == 18)
||(x_pointer == 53 && y_pointer == 18)
||(x_pointer == 54 && y_pointer == 18)
||(x_pointer == 55 && y_pointer == 18)
||(x_pointer == 56 && y_pointer == 18)
||(x_pointer == 57 && y_pointer == 18)
||(x_pointer == 58 && y_pointer == 18)
||(x_pointer == 68 && y_pointer == 18)
||(x_pointer == 69 && y_pointer == 18)
||(x_pointer == 70 && y_pointer == 18)
||(x_pointer == 71 && y_pointer == 18)
||(x_pointer == 72 && y_pointer == 18)
||(x_pointer == 73 && y_pointer == 18)
||(x_pointer == 74 && y_pointer == 18)
||(x_pointer == 75 && y_pointer == 18)
||(x_pointer == 76 && y_pointer == 18)
||(x_pointer == 77 && y_pointer == 18)
||(x_pointer == 78 && y_pointer == 18)
||(x_pointer == 79 && y_pointer == 18)
||(x_pointer == 80 && y_pointer == 18)
||(x_pointer == 81 && y_pointer == 18)
||(x_pointer == 82 && y_pointer == 18)
||(x_pointer == 83 && y_pointer == 18)
||(x_pointer == 84 && y_pointer == 18)
||(x_pointer == 85 && y_pointer == 18)
||(x_pointer == 86 && y_pointer == 18)
||(x_pointer == 87 && y_pointer == 18)
||(x_pointer == 88 && y_pointer == 18)
||(x_pointer == 89 && y_pointer == 18)
||(x_pointer == 90 && y_pointer == 18)
||(x_pointer == 91 && y_pointer == 18)
||(x_pointer == 92 && y_pointer == 18)
||(x_pointer == 93 && y_pointer == 18)
||(x_pointer == 94 && y_pointer == 18)
||(x_pointer == 95 && y_pointer == 18)
||(x_pointer == 96 && y_pointer == 18)
||(x_pointer == 97 && y_pointer == 18)
||(x_pointer == 98 && y_pointer == 18)
||(x_pointer == 99 && y_pointer == 18)
||(x_pointer == 100 && y_pointer == 18)
||(x_pointer == 101 && y_pointer == 18)
||(x_pointer == 102 && y_pointer == 18)
||(x_pointer == 103 && y_pointer == 18)
||(x_pointer == 104 && y_pointer == 18)
||(x_pointer == 105 && y_pointer == 18)
||(x_pointer == 106 && y_pointer == 18)
||(x_pointer == 107 && y_pointer == 18)
||(x_pointer == 108 && y_pointer == 18)
||(x_pointer == 109 && y_pointer == 18)
||(x_pointer == 110 && y_pointer == 18)
||(x_pointer == 111 && y_pointer == 18)
||(x_pointer == 112 && y_pointer == 18)
||(x_pointer == 113 && y_pointer == 18)
||(x_pointer == 114 && y_pointer == 18)
||(x_pointer == 115 && y_pointer == 18)
||(x_pointer == 116 && y_pointer == 18)
||(x_pointer == 117 && y_pointer == 18)
||(x_pointer == 118 && y_pointer == 18)
||(x_pointer == 119 && y_pointer == 18)
||(x_pointer == 120 && y_pointer == 18)
||(x_pointer == 121 && y_pointer == 18)
||(x_pointer == 122 && y_pointer == 18)
||(x_pointer == 123 && y_pointer == 18)
||(x_pointer == 124 && y_pointer == 18)
||(x_pointer == 125 && y_pointer == 18)
||(x_pointer == 126 && y_pointer == 18)
||(x_pointer == 127 && y_pointer == 18)
||(x_pointer == 128 && y_pointer == 18)
||(x_pointer == 129 && y_pointer == 18)
||(x_pointer == 130 && y_pointer == 18)
||(x_pointer == 131 && y_pointer == 18)
||(x_pointer == 132 && y_pointer == 18)
||(x_pointer == 133 && y_pointer == 18)
||(x_pointer == 134 && y_pointer == 18)
||(x_pointer == 135 && y_pointer == 18)
||(x_pointer == 136 && y_pointer == 18)
||(x_pointer == 137 && y_pointer == 18)
||(x_pointer == 138 && y_pointer == 18)
||(x_pointer == 139 && y_pointer == 18)
||(x_pointer == 140 && y_pointer == 18)
||(x_pointer == 141 && y_pointer == 18)
||(x_pointer == 142 && y_pointer == 18)
||(x_pointer == 143 && y_pointer == 18)
||(x_pointer == 144 && y_pointer == 18)
||(x_pointer == 145 && y_pointer == 18)
||(x_pointer == 14 && y_pointer == 19)
||(x_pointer == 15 && y_pointer == 19)
||(x_pointer == 16 && y_pointer == 19)
||(x_pointer == 26 && y_pointer == 19)
||(x_pointer == 27 && y_pointer == 19)
||(x_pointer == 28 && y_pointer == 19)
||(x_pointer == 29 && y_pointer == 19)
||(x_pointer == 30 && y_pointer == 19)
||(x_pointer == 31 && y_pointer == 19)
||(x_pointer == 32 && y_pointer == 19)
||(x_pointer == 33 && y_pointer == 19)
||(x_pointer == 34 && y_pointer == 19)
||(x_pointer == 35 && y_pointer == 19)
||(x_pointer == 36 && y_pointer == 19)
||(x_pointer == 37 && y_pointer == 19)
||(x_pointer == 38 && y_pointer == 19)
||(x_pointer == 39 && y_pointer == 19)
||(x_pointer == 40 && y_pointer == 19)
||(x_pointer == 41 && y_pointer == 19)
||(x_pointer == 42 && y_pointer == 19)
||(x_pointer == 43 && y_pointer == 19)
||(x_pointer == 53 && y_pointer == 19)
||(x_pointer == 54 && y_pointer == 19)
||(x_pointer == 55 && y_pointer == 19)
||(x_pointer == 56 && y_pointer == 19)
||(x_pointer == 57 && y_pointer == 19)
||(x_pointer == 58 && y_pointer == 19)
||(x_pointer == 68 && y_pointer == 19)
||(x_pointer == 69 && y_pointer == 19)
||(x_pointer == 70 && y_pointer == 19)
||(x_pointer == 71 && y_pointer == 19)
||(x_pointer == 72 && y_pointer == 19)
||(x_pointer == 73 && y_pointer == 19)
||(x_pointer == 74 && y_pointer == 19)
||(x_pointer == 75 && y_pointer == 19)
||(x_pointer == 76 && y_pointer == 19)
||(x_pointer == 77 && y_pointer == 19)
||(x_pointer == 78 && y_pointer == 19)
||(x_pointer == 79 && y_pointer == 19)
||(x_pointer == 80 && y_pointer == 19)
||(x_pointer == 81 && y_pointer == 19)
||(x_pointer == 82 && y_pointer == 19)
||(x_pointer == 83 && y_pointer == 19)
||(x_pointer == 84 && y_pointer == 19)
||(x_pointer == 85 && y_pointer == 19)
||(x_pointer == 86 && y_pointer == 19)
||(x_pointer == 87 && y_pointer == 19)
||(x_pointer == 88 && y_pointer == 19)
||(x_pointer == 89 && y_pointer == 19)
||(x_pointer == 90 && y_pointer == 19)
||(x_pointer == 91 && y_pointer == 19)
||(x_pointer == 92 && y_pointer == 19)
||(x_pointer == 93 && y_pointer == 19)
||(x_pointer == 94 && y_pointer == 19)
||(x_pointer == 95 && y_pointer == 19)
||(x_pointer == 96 && y_pointer == 19)
||(x_pointer == 97 && y_pointer == 19)
||(x_pointer == 98 && y_pointer == 19)
||(x_pointer == 99 && y_pointer == 19)
||(x_pointer == 100 && y_pointer == 19)
||(x_pointer == 101 && y_pointer == 19)
||(x_pointer == 102 && y_pointer == 19)
||(x_pointer == 103 && y_pointer == 19)
||(x_pointer == 104 && y_pointer == 19)
||(x_pointer == 105 && y_pointer == 19)
||(x_pointer == 106 && y_pointer == 19)
||(x_pointer == 107 && y_pointer == 19)
||(x_pointer == 108 && y_pointer == 19)
||(x_pointer == 109 && y_pointer == 19)
||(x_pointer == 110 && y_pointer == 19)
||(x_pointer == 111 && y_pointer == 19)
||(x_pointer == 112 && y_pointer == 19)
||(x_pointer == 113 && y_pointer == 19)
||(x_pointer == 114 && y_pointer == 19)
||(x_pointer == 115 && y_pointer == 19)
||(x_pointer == 116 && y_pointer == 19)
||(x_pointer == 117 && y_pointer == 19)
||(x_pointer == 118 && y_pointer == 19)
||(x_pointer == 119 && y_pointer == 19)
||(x_pointer == 120 && y_pointer == 19)
||(x_pointer == 121 && y_pointer == 19)
||(x_pointer == 122 && y_pointer == 19)
||(x_pointer == 123 && y_pointer == 19)
||(x_pointer == 124 && y_pointer == 19)
||(x_pointer == 125 && y_pointer == 19)
||(x_pointer == 126 && y_pointer == 19)
||(x_pointer == 127 && y_pointer == 19)
||(x_pointer == 128 && y_pointer == 19)
||(x_pointer == 129 && y_pointer == 19)
||(x_pointer == 130 && y_pointer == 19)
||(x_pointer == 131 && y_pointer == 19)
||(x_pointer == 132 && y_pointer == 19)
||(x_pointer == 133 && y_pointer == 19)
||(x_pointer == 134 && y_pointer == 19)
||(x_pointer == 135 && y_pointer == 19)
||(x_pointer == 136 && y_pointer == 19)
||(x_pointer == 137 && y_pointer == 19)
||(x_pointer == 138 && y_pointer == 19)
||(x_pointer == 139 && y_pointer == 19)
||(x_pointer == 140 && y_pointer == 19)
||(x_pointer == 141 && y_pointer == 19)
||(x_pointer == 142 && y_pointer == 19)
||(x_pointer == 143 && y_pointer == 19)
||(x_pointer == 144 && y_pointer == 19)
||(x_pointer == 145 && y_pointer == 19)
||(x_pointer == 14 && y_pointer == 20)
||(x_pointer == 15 && y_pointer == 20)
||(x_pointer == 16 && y_pointer == 20)
||(x_pointer == 26 && y_pointer == 20)
||(x_pointer == 27 && y_pointer == 20)
||(x_pointer == 28 && y_pointer == 20)
||(x_pointer == 56 && y_pointer == 20)
||(x_pointer == 57 && y_pointer == 20)
||(x_pointer == 58 && y_pointer == 20)
||(x_pointer == 68 && y_pointer == 20)
||(x_pointer == 69 && y_pointer == 20)
||(x_pointer == 70 && y_pointer == 20)
||(x_pointer == 143 && y_pointer == 20)
||(x_pointer == 144 && y_pointer == 20)
||(x_pointer == 145 && y_pointer == 20)
||(x_pointer == 14 && y_pointer == 21)
||(x_pointer == 15 && y_pointer == 21)
||(x_pointer == 16 && y_pointer == 21)
||(x_pointer == 26 && y_pointer == 21)
||(x_pointer == 27 && y_pointer == 21)
||(x_pointer == 28 && y_pointer == 21)
||(x_pointer == 56 && y_pointer == 21)
||(x_pointer == 57 && y_pointer == 21)
||(x_pointer == 58 && y_pointer == 21)
||(x_pointer == 68 && y_pointer == 21)
||(x_pointer == 69 && y_pointer == 21)
||(x_pointer == 70 && y_pointer == 21)
||(x_pointer == 143 && y_pointer == 21)
||(x_pointer == 144 && y_pointer == 21)
||(x_pointer == 145 && y_pointer == 21)
||(x_pointer == 14 && y_pointer == 22)
||(x_pointer == 15 && y_pointer == 22)
||(x_pointer == 16 && y_pointer == 22)
||(x_pointer == 26 && y_pointer == 22)
||(x_pointer == 27 && y_pointer == 22)
||(x_pointer == 28 && y_pointer == 22)
||(x_pointer == 56 && y_pointer == 22)
||(x_pointer == 57 && y_pointer == 22)
||(x_pointer == 58 && y_pointer == 22)
||(x_pointer == 68 && y_pointer == 22)
||(x_pointer == 69 && y_pointer == 22)
||(x_pointer == 70 && y_pointer == 22)
||(x_pointer == 143 && y_pointer == 22)
||(x_pointer == 144 && y_pointer == 22)
||(x_pointer == 145 && y_pointer == 22)
||(x_pointer == 14 && y_pointer == 23)
||(x_pointer == 15 && y_pointer == 23)
||(x_pointer == 16 && y_pointer == 23)
||(x_pointer == 26 && y_pointer == 23)
||(x_pointer == 27 && y_pointer == 23)
||(x_pointer == 28 && y_pointer == 23)
||(x_pointer == 56 && y_pointer == 23)
||(x_pointer == 57 && y_pointer == 23)
||(x_pointer == 58 && y_pointer == 23)
||(x_pointer == 68 && y_pointer == 23)
||(x_pointer == 69 && y_pointer == 23)
||(x_pointer == 70 && y_pointer == 23)
||(x_pointer == 143 && y_pointer == 23)
||(x_pointer == 144 && y_pointer == 23)
||(x_pointer == 145 && y_pointer == 23)
||(x_pointer == 14 && y_pointer == 24)
||(x_pointer == 15 && y_pointer == 24)
||(x_pointer == 16 && y_pointer == 24)
||(x_pointer == 26 && y_pointer == 24)
||(x_pointer == 27 && y_pointer == 24)
||(x_pointer == 28 && y_pointer == 24)
||(x_pointer == 56 && y_pointer == 24)
||(x_pointer == 57 && y_pointer == 24)
||(x_pointer == 58 && y_pointer == 24)
||(x_pointer == 68 && y_pointer == 24)
||(x_pointer == 69 && y_pointer == 24)
||(x_pointer == 70 && y_pointer == 24)
||(x_pointer == 143 && y_pointer == 24)
||(x_pointer == 144 && y_pointer == 24)
||(x_pointer == 145 && y_pointer == 24)
||(x_pointer == 14 && y_pointer == 25)
||(x_pointer == 15 && y_pointer == 25)
||(x_pointer == 16 && y_pointer == 25)
||(x_pointer == 26 && y_pointer == 25)
||(x_pointer == 27 && y_pointer == 25)
||(x_pointer == 28 && y_pointer == 25)
||(x_pointer == 56 && y_pointer == 25)
||(x_pointer == 57 && y_pointer == 25)
||(x_pointer == 58 && y_pointer == 25)
||(x_pointer == 68 && y_pointer == 25)
||(x_pointer == 69 && y_pointer == 25)
||(x_pointer == 70 && y_pointer == 25)
||(x_pointer == 143 && y_pointer == 25)
||(x_pointer == 144 && y_pointer == 25)
||(x_pointer == 145 && y_pointer == 25)
||(x_pointer == 14 && y_pointer == 26)
||(x_pointer == 15 && y_pointer == 26)
||(x_pointer == 16 && y_pointer == 26)
||(x_pointer == 53 && y_pointer == 26)
||(x_pointer == 54 && y_pointer == 26)
||(x_pointer == 55 && y_pointer == 26)
||(x_pointer == 56 && y_pointer == 26)
||(x_pointer == 57 && y_pointer == 26)
||(x_pointer == 58 && y_pointer == 26)
||(x_pointer == 68 && y_pointer == 26)
||(x_pointer == 69 && y_pointer == 26)
||(x_pointer == 70 && y_pointer == 26)
||(x_pointer == 143 && y_pointer == 26)
||(x_pointer == 144 && y_pointer == 26)
||(x_pointer == 145 && y_pointer == 26)
||(x_pointer == 14 && y_pointer == 27)
||(x_pointer == 15 && y_pointer == 27)
||(x_pointer == 16 && y_pointer == 27)
||(x_pointer == 53 && y_pointer == 27)
||(x_pointer == 54 && y_pointer == 27)
||(x_pointer == 55 && y_pointer == 27)
||(x_pointer == 56 && y_pointer == 27)
||(x_pointer == 57 && y_pointer == 27)
||(x_pointer == 58 && y_pointer == 27)
||(x_pointer == 68 && y_pointer == 27)
||(x_pointer == 69 && y_pointer == 27)
||(x_pointer == 70 && y_pointer == 27)
||(x_pointer == 143 && y_pointer == 27)
||(x_pointer == 144 && y_pointer == 27)
||(x_pointer == 145 && y_pointer == 27)
||(x_pointer == 14 && y_pointer == 28)
||(x_pointer == 15 && y_pointer == 28)
||(x_pointer == 16 && y_pointer == 28)
||(x_pointer == 53 && y_pointer == 28)
||(x_pointer == 54 && y_pointer == 28)
||(x_pointer == 55 && y_pointer == 28)
||(x_pointer == 56 && y_pointer == 28)
||(x_pointer == 57 && y_pointer == 28)
||(x_pointer == 58 && y_pointer == 28)
||(x_pointer == 68 && y_pointer == 28)
||(x_pointer == 69 && y_pointer == 28)
||(x_pointer == 70 && y_pointer == 28)
||(x_pointer == 143 && y_pointer == 28)
||(x_pointer == 144 && y_pointer == 28)
||(x_pointer == 145 && y_pointer == 28)
||(x_pointer == 14 && y_pointer == 29)
||(x_pointer == 15 && y_pointer == 29)
||(x_pointer == 16 && y_pointer == 29)
||(x_pointer == 68 && y_pointer == 29)
||(x_pointer == 69 && y_pointer == 29)
||(x_pointer == 70 && y_pointer == 29)
||(x_pointer == 83 && y_pointer == 29)
||(x_pointer == 84 && y_pointer == 29)
||(x_pointer == 85 && y_pointer == 29)
||(x_pointer == 86 && y_pointer == 29)
||(x_pointer == 87 && y_pointer == 29)
||(x_pointer == 88 && y_pointer == 29)
||(x_pointer == 89 && y_pointer == 29)
||(x_pointer == 90 && y_pointer == 29)
||(x_pointer == 91 && y_pointer == 29)
||(x_pointer == 92 && y_pointer == 29)
||(x_pointer == 93 && y_pointer == 29)
||(x_pointer == 94 && y_pointer == 29)
||(x_pointer == 95 && y_pointer == 29)
||(x_pointer == 96 && y_pointer == 29)
||(x_pointer == 97 && y_pointer == 29)
||(x_pointer == 98 && y_pointer == 29)
||(x_pointer == 99 && y_pointer == 29)
||(x_pointer == 100 && y_pointer == 29)
||(x_pointer == 101 && y_pointer == 29)
||(x_pointer == 102 && y_pointer == 29)
||(x_pointer == 103 && y_pointer == 29)
||(x_pointer == 104 && y_pointer == 29)
||(x_pointer == 105 && y_pointer == 29)
||(x_pointer == 106 && y_pointer == 29)
||(x_pointer == 107 && y_pointer == 29)
||(x_pointer == 108 && y_pointer == 29)
||(x_pointer == 109 && y_pointer == 29)
||(x_pointer == 110 && y_pointer == 29)
||(x_pointer == 111 && y_pointer == 29)
||(x_pointer == 112 && y_pointer == 29)
||(x_pointer == 113 && y_pointer == 29)
||(x_pointer == 114 && y_pointer == 29)
||(x_pointer == 115 && y_pointer == 29)
||(x_pointer == 116 && y_pointer == 29)
||(x_pointer == 117 && y_pointer == 29)
||(x_pointer == 118 && y_pointer == 29)
||(x_pointer == 119 && y_pointer == 29)
||(x_pointer == 120 && y_pointer == 29)
||(x_pointer == 121 && y_pointer == 29)
||(x_pointer == 122 && y_pointer == 29)
||(x_pointer == 123 && y_pointer == 29)
||(x_pointer == 124 && y_pointer == 29)
||(x_pointer == 125 && y_pointer == 29)
||(x_pointer == 126 && y_pointer == 29)
||(x_pointer == 127 && y_pointer == 29)
||(x_pointer == 128 && y_pointer == 29)
||(x_pointer == 129 && y_pointer == 29)
||(x_pointer == 130 && y_pointer == 29)
||(x_pointer == 131 && y_pointer == 29)
||(x_pointer == 132 && y_pointer == 29)
||(x_pointer == 133 && y_pointer == 29)
||(x_pointer == 134 && y_pointer == 29)
||(x_pointer == 135 && y_pointer == 29)
||(x_pointer == 136 && y_pointer == 29)
||(x_pointer == 137 && y_pointer == 29)
||(x_pointer == 138 && y_pointer == 29)
||(x_pointer == 139 && y_pointer == 29)
||(x_pointer == 140 && y_pointer == 29)
||(x_pointer == 141 && y_pointer == 29)
||(x_pointer == 142 && y_pointer == 29)
||(x_pointer == 143 && y_pointer == 29)
||(x_pointer == 144 && y_pointer == 29)
||(x_pointer == 145 && y_pointer == 29)
||(x_pointer == 14 && y_pointer == 30)
||(x_pointer == 15 && y_pointer == 30)
||(x_pointer == 16 && y_pointer == 30)
||(x_pointer == 68 && y_pointer == 30)
||(x_pointer == 69 && y_pointer == 30)
||(x_pointer == 70 && y_pointer == 30)
||(x_pointer == 83 && y_pointer == 30)
||(x_pointer == 84 && y_pointer == 30)
||(x_pointer == 85 && y_pointer == 30)
||(x_pointer == 86 && y_pointer == 30)
||(x_pointer == 87 && y_pointer == 30)
||(x_pointer == 88 && y_pointer == 30)
||(x_pointer == 89 && y_pointer == 30)
||(x_pointer == 90 && y_pointer == 30)
||(x_pointer == 91 && y_pointer == 30)
||(x_pointer == 92 && y_pointer == 30)
||(x_pointer == 93 && y_pointer == 30)
||(x_pointer == 94 && y_pointer == 30)
||(x_pointer == 95 && y_pointer == 30)
||(x_pointer == 96 && y_pointer == 30)
||(x_pointer == 97 && y_pointer == 30)
||(x_pointer == 98 && y_pointer == 30)
||(x_pointer == 99 && y_pointer == 30)
||(x_pointer == 100 && y_pointer == 30)
||(x_pointer == 101 && y_pointer == 30)
||(x_pointer == 102 && y_pointer == 30)
||(x_pointer == 103 && y_pointer == 30)
||(x_pointer == 104 && y_pointer == 30)
||(x_pointer == 105 && y_pointer == 30)
||(x_pointer == 106 && y_pointer == 30)
||(x_pointer == 107 && y_pointer == 30)
||(x_pointer == 108 && y_pointer == 30)
||(x_pointer == 109 && y_pointer == 30)
||(x_pointer == 110 && y_pointer == 30)
||(x_pointer == 111 && y_pointer == 30)
||(x_pointer == 112 && y_pointer == 30)
||(x_pointer == 113 && y_pointer == 30)
||(x_pointer == 114 && y_pointer == 30)
||(x_pointer == 115 && y_pointer == 30)
||(x_pointer == 116 && y_pointer == 30)
||(x_pointer == 117 && y_pointer == 30)
||(x_pointer == 118 && y_pointer == 30)
||(x_pointer == 119 && y_pointer == 30)
||(x_pointer == 120 && y_pointer == 30)
||(x_pointer == 121 && y_pointer == 30)
||(x_pointer == 122 && y_pointer == 30)
||(x_pointer == 123 && y_pointer == 30)
||(x_pointer == 124 && y_pointer == 30)
||(x_pointer == 125 && y_pointer == 30)
||(x_pointer == 126 && y_pointer == 30)
||(x_pointer == 127 && y_pointer == 30)
||(x_pointer == 128 && y_pointer == 30)
||(x_pointer == 129 && y_pointer == 30)
||(x_pointer == 130 && y_pointer == 30)
||(x_pointer == 131 && y_pointer == 30)
||(x_pointer == 132 && y_pointer == 30)
||(x_pointer == 133 && y_pointer == 30)
||(x_pointer == 134 && y_pointer == 30)
||(x_pointer == 135 && y_pointer == 30)
||(x_pointer == 136 && y_pointer == 30)
||(x_pointer == 137 && y_pointer == 30)
||(x_pointer == 138 && y_pointer == 30)
||(x_pointer == 139 && y_pointer == 30)
||(x_pointer == 140 && y_pointer == 30)
||(x_pointer == 141 && y_pointer == 30)
||(x_pointer == 142 && y_pointer == 30)
||(x_pointer == 143 && y_pointer == 30)
||(x_pointer == 144 && y_pointer == 30)
||(x_pointer == 145 && y_pointer == 30)
||(x_pointer == 14 && y_pointer == 31)
||(x_pointer == 15 && y_pointer == 31)
||(x_pointer == 16 && y_pointer == 31)
||(x_pointer == 68 && y_pointer == 31)
||(x_pointer == 69 && y_pointer == 31)
||(x_pointer == 70 && y_pointer == 31)
||(x_pointer == 83 && y_pointer == 31)
||(x_pointer == 84 && y_pointer == 31)
||(x_pointer == 85 && y_pointer == 31)
||(x_pointer == 86 && y_pointer == 31)
||(x_pointer == 87 && y_pointer == 31)
||(x_pointer == 88 && y_pointer == 31)
||(x_pointer == 89 && y_pointer == 31)
||(x_pointer == 90 && y_pointer == 31)
||(x_pointer == 91 && y_pointer == 31)
||(x_pointer == 92 && y_pointer == 31)
||(x_pointer == 93 && y_pointer == 31)
||(x_pointer == 94 && y_pointer == 31)
||(x_pointer == 95 && y_pointer == 31)
||(x_pointer == 96 && y_pointer == 31)
||(x_pointer == 97 && y_pointer == 31)
||(x_pointer == 98 && y_pointer == 31)
||(x_pointer == 99 && y_pointer == 31)
||(x_pointer == 100 && y_pointer == 31)
||(x_pointer == 101 && y_pointer == 31)
||(x_pointer == 102 && y_pointer == 31)
||(x_pointer == 103 && y_pointer == 31)
||(x_pointer == 104 && y_pointer == 31)
||(x_pointer == 105 && y_pointer == 31)
||(x_pointer == 106 && y_pointer == 31)
||(x_pointer == 107 && y_pointer == 31)
||(x_pointer == 108 && y_pointer == 31)
||(x_pointer == 109 && y_pointer == 31)
||(x_pointer == 110 && y_pointer == 31)
||(x_pointer == 111 && y_pointer == 31)
||(x_pointer == 112 && y_pointer == 31)
||(x_pointer == 113 && y_pointer == 31)
||(x_pointer == 114 && y_pointer == 31)
||(x_pointer == 115 && y_pointer == 31)
||(x_pointer == 116 && y_pointer == 31)
||(x_pointer == 117 && y_pointer == 31)
||(x_pointer == 118 && y_pointer == 31)
||(x_pointer == 119 && y_pointer == 31)
||(x_pointer == 120 && y_pointer == 31)
||(x_pointer == 121 && y_pointer == 31)
||(x_pointer == 122 && y_pointer == 31)
||(x_pointer == 123 && y_pointer == 31)
||(x_pointer == 124 && y_pointer == 31)
||(x_pointer == 125 && y_pointer == 31)
||(x_pointer == 126 && y_pointer == 31)
||(x_pointer == 127 && y_pointer == 31)
||(x_pointer == 128 && y_pointer == 31)
||(x_pointer == 129 && y_pointer == 31)
||(x_pointer == 130 && y_pointer == 31)
||(x_pointer == 131 && y_pointer == 31)
||(x_pointer == 132 && y_pointer == 31)
||(x_pointer == 133 && y_pointer == 31)
||(x_pointer == 134 && y_pointer == 31)
||(x_pointer == 135 && y_pointer == 31)
||(x_pointer == 136 && y_pointer == 31)
||(x_pointer == 137 && y_pointer == 31)
||(x_pointer == 138 && y_pointer == 31)
||(x_pointer == 139 && y_pointer == 31)
||(x_pointer == 140 && y_pointer == 31)
||(x_pointer == 141 && y_pointer == 31)
||(x_pointer == 142 && y_pointer == 31)
||(x_pointer == 143 && y_pointer == 31)
||(x_pointer == 144 && y_pointer == 31)
||(x_pointer == 145 && y_pointer == 31)
||(x_pointer == 14 && y_pointer == 32)
||(x_pointer == 15 && y_pointer == 32)
||(x_pointer == 16 && y_pointer == 32)
||(x_pointer == 68 && y_pointer == 32)
||(x_pointer == 69 && y_pointer == 32)
||(x_pointer == 70 && y_pointer == 32)
||(x_pointer == 83 && y_pointer == 32)
||(x_pointer == 84 && y_pointer == 32)
||(x_pointer == 85 && y_pointer == 32)
||(x_pointer == 14 && y_pointer == 33)
||(x_pointer == 15 && y_pointer == 33)
||(x_pointer == 16 && y_pointer == 33)
||(x_pointer == 68 && y_pointer == 33)
||(x_pointer == 69 && y_pointer == 33)
||(x_pointer == 70 && y_pointer == 33)
||(x_pointer == 83 && y_pointer == 33)
||(x_pointer == 84 && y_pointer == 33)
||(x_pointer == 85 && y_pointer == 33)
||(x_pointer == 14 && y_pointer == 34)
||(x_pointer == 15 && y_pointer == 34)
||(x_pointer == 16 && y_pointer == 34)
||(x_pointer == 68 && y_pointer == 34)
||(x_pointer == 69 && y_pointer == 34)
||(x_pointer == 70 && y_pointer == 34)
||(x_pointer == 83 && y_pointer == 34)
||(x_pointer == 84 && y_pointer == 34)
||(x_pointer == 85 && y_pointer == 34)
||(x_pointer == 14 && y_pointer == 35)
||(x_pointer == 15 && y_pointer == 35)
||(x_pointer == 16 && y_pointer == 35)
||(x_pointer == 68 && y_pointer == 35)
||(x_pointer == 69 && y_pointer == 35)
||(x_pointer == 70 && y_pointer == 35)
||(x_pointer == 83 && y_pointer == 35)
||(x_pointer == 84 && y_pointer == 35)
||(x_pointer == 85 && y_pointer == 35)
||(x_pointer == 14 && y_pointer == 36)
||(x_pointer == 15 && y_pointer == 36)
||(x_pointer == 16 && y_pointer == 36)
||(x_pointer == 68 && y_pointer == 36)
||(x_pointer == 69 && y_pointer == 36)
||(x_pointer == 70 && y_pointer == 36)
||(x_pointer == 83 && y_pointer == 36)
||(x_pointer == 84 && y_pointer == 36)
||(x_pointer == 85 && y_pointer == 36)
||(x_pointer == 14 && y_pointer == 37)
||(x_pointer == 15 && y_pointer == 37)
||(x_pointer == 16 && y_pointer == 37)
||(x_pointer == 68 && y_pointer == 37)
||(x_pointer == 69 && y_pointer == 37)
||(x_pointer == 70 && y_pointer == 37)
||(x_pointer == 83 && y_pointer == 37)
||(x_pointer == 84 && y_pointer == 37)
||(x_pointer == 85 && y_pointer == 37)
||(x_pointer == 14 && y_pointer == 38)
||(x_pointer == 15 && y_pointer == 38)
||(x_pointer == 16 && y_pointer == 38)
||(x_pointer == 53 && y_pointer == 38)
||(x_pointer == 54 && y_pointer == 38)
||(x_pointer == 55 && y_pointer == 38)
||(x_pointer == 56 && y_pointer == 38)
||(x_pointer == 57 && y_pointer == 38)
||(x_pointer == 58 && y_pointer == 38)
||(x_pointer == 59 && y_pointer == 38)
||(x_pointer == 60 && y_pointer == 38)
||(x_pointer == 61 && y_pointer == 38)
||(x_pointer == 62 && y_pointer == 38)
||(x_pointer == 63 && y_pointer == 38)
||(x_pointer == 64 && y_pointer == 38)
||(x_pointer == 65 && y_pointer == 38)
||(x_pointer == 66 && y_pointer == 38)
||(x_pointer == 67 && y_pointer == 38)
||(x_pointer == 68 && y_pointer == 38)
||(x_pointer == 69 && y_pointer == 38)
||(x_pointer == 70 && y_pointer == 38)
||(x_pointer == 83 && y_pointer == 38)
||(x_pointer == 84 && y_pointer == 38)
||(x_pointer == 85 && y_pointer == 38)
||(x_pointer == 14 && y_pointer == 39)
||(x_pointer == 15 && y_pointer == 39)
||(x_pointer == 16 && y_pointer == 39)
||(x_pointer == 53 && y_pointer == 39)
||(x_pointer == 54 && y_pointer == 39)
||(x_pointer == 55 && y_pointer == 39)
||(x_pointer == 56 && y_pointer == 39)
||(x_pointer == 57 && y_pointer == 39)
||(x_pointer == 58 && y_pointer == 39)
||(x_pointer == 59 && y_pointer == 39)
||(x_pointer == 60 && y_pointer == 39)
||(x_pointer == 61 && y_pointer == 39)
||(x_pointer == 62 && y_pointer == 39)
||(x_pointer == 63 && y_pointer == 39)
||(x_pointer == 64 && y_pointer == 39)
||(x_pointer == 65 && y_pointer == 39)
||(x_pointer == 66 && y_pointer == 39)
||(x_pointer == 67 && y_pointer == 39)
||(x_pointer == 68 && y_pointer == 39)
||(x_pointer == 69 && y_pointer == 39)
||(x_pointer == 70 && y_pointer == 39)
||(x_pointer == 83 && y_pointer == 39)
||(x_pointer == 84 && y_pointer == 39)
||(x_pointer == 85 && y_pointer == 39)
||(x_pointer == 14 && y_pointer == 40)
||(x_pointer == 15 && y_pointer == 40)
||(x_pointer == 16 && y_pointer == 40)
||(x_pointer == 53 && y_pointer == 40)
||(x_pointer == 54 && y_pointer == 40)
||(x_pointer == 55 && y_pointer == 40)
||(x_pointer == 56 && y_pointer == 40)
||(x_pointer == 57 && y_pointer == 40)
||(x_pointer == 58 && y_pointer == 40)
||(x_pointer == 59 && y_pointer == 40)
||(x_pointer == 60 && y_pointer == 40)
||(x_pointer == 61 && y_pointer == 40)
||(x_pointer == 62 && y_pointer == 40)
||(x_pointer == 63 && y_pointer == 40)
||(x_pointer == 64 && y_pointer == 40)
||(x_pointer == 65 && y_pointer == 40)
||(x_pointer == 66 && y_pointer == 40)
||(x_pointer == 67 && y_pointer == 40)
||(x_pointer == 68 && y_pointer == 40)
||(x_pointer == 69 && y_pointer == 40)
||(x_pointer == 70 && y_pointer == 40)
||(x_pointer == 83 && y_pointer == 40)
||(x_pointer == 84 && y_pointer == 40)
||(x_pointer == 85 && y_pointer == 40)
||(x_pointer == 14 && y_pointer == 41)
||(x_pointer == 15 && y_pointer == 41)
||(x_pointer == 16 && y_pointer == 41)
||(x_pointer == 26 && y_pointer == 41)
||(x_pointer == 27 && y_pointer == 41)
||(x_pointer == 28 && y_pointer == 41)
||(x_pointer == 95 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 99 && y_pointer == 41)
||(x_pointer == 100 && y_pointer == 41)
||(x_pointer == 101 && y_pointer == 41)
||(x_pointer == 102 && y_pointer == 41)
||(x_pointer == 103 && y_pointer == 41)
||(x_pointer == 104 && y_pointer == 41)
||(x_pointer == 105 && y_pointer == 41)
||(x_pointer == 106 && y_pointer == 41)
||(x_pointer == 107 && y_pointer == 41)
||(x_pointer == 108 && y_pointer == 41)
||(x_pointer == 109 && y_pointer == 41)
||(x_pointer == 110 && y_pointer == 41)
||(x_pointer == 111 && y_pointer == 41)
||(x_pointer == 112 && y_pointer == 41)
||(x_pointer == 113 && y_pointer == 41)
||(x_pointer == 114 && y_pointer == 41)
||(x_pointer == 115 && y_pointer == 41)
||(x_pointer == 116 && y_pointer == 41)
||(x_pointer == 117 && y_pointer == 41)
||(x_pointer == 118 && y_pointer == 41)
||(x_pointer == 119 && y_pointer == 41)
||(x_pointer == 120 && y_pointer == 41)
||(x_pointer == 121 && y_pointer == 41)
||(x_pointer == 122 && y_pointer == 41)
||(x_pointer == 123 && y_pointer == 41)
||(x_pointer == 124 && y_pointer == 41)
||(x_pointer == 125 && y_pointer == 41)
||(x_pointer == 126 && y_pointer == 41)
||(x_pointer == 127 && y_pointer == 41)
||(x_pointer == 128 && y_pointer == 41)
||(x_pointer == 129 && y_pointer == 41)
||(x_pointer == 130 && y_pointer == 41)
||(x_pointer == 131 && y_pointer == 41)
||(x_pointer == 132 && y_pointer == 41)
||(x_pointer == 133 && y_pointer == 41)
||(x_pointer == 134 && y_pointer == 41)
||(x_pointer == 135 && y_pointer == 41)
||(x_pointer == 136 && y_pointer == 41)
||(x_pointer == 137 && y_pointer == 41)
||(x_pointer == 138 && y_pointer == 41)
||(x_pointer == 139 && y_pointer == 41)
||(x_pointer == 140 && y_pointer == 41)
||(x_pointer == 141 && y_pointer == 41)
||(x_pointer == 142 && y_pointer == 41)
||(x_pointer == 143 && y_pointer == 41)
||(x_pointer == 144 && y_pointer == 41)
||(x_pointer == 145 && y_pointer == 41)
||(x_pointer == 14 && y_pointer == 42)
||(x_pointer == 15 && y_pointer == 42)
||(x_pointer == 16 && y_pointer == 42)
||(x_pointer == 26 && y_pointer == 42)
||(x_pointer == 27 && y_pointer == 42)
||(x_pointer == 28 && y_pointer == 42)
||(x_pointer == 95 && y_pointer == 42)
||(x_pointer == 96 && y_pointer == 42)
||(x_pointer == 97 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 99 && y_pointer == 42)
||(x_pointer == 100 && y_pointer == 42)
||(x_pointer == 101 && y_pointer == 42)
||(x_pointer == 102 && y_pointer == 42)
||(x_pointer == 103 && y_pointer == 42)
||(x_pointer == 104 && y_pointer == 42)
||(x_pointer == 105 && y_pointer == 42)
||(x_pointer == 106 && y_pointer == 42)
||(x_pointer == 107 && y_pointer == 42)
||(x_pointer == 108 && y_pointer == 42)
||(x_pointer == 109 && y_pointer == 42)
||(x_pointer == 110 && y_pointer == 42)
||(x_pointer == 111 && y_pointer == 42)
||(x_pointer == 112 && y_pointer == 42)
||(x_pointer == 113 && y_pointer == 42)
||(x_pointer == 114 && y_pointer == 42)
||(x_pointer == 115 && y_pointer == 42)
||(x_pointer == 116 && y_pointer == 42)
||(x_pointer == 117 && y_pointer == 42)
||(x_pointer == 118 && y_pointer == 42)
||(x_pointer == 119 && y_pointer == 42)
||(x_pointer == 120 && y_pointer == 42)
||(x_pointer == 121 && y_pointer == 42)
||(x_pointer == 122 && y_pointer == 42)
||(x_pointer == 123 && y_pointer == 42)
||(x_pointer == 124 && y_pointer == 42)
||(x_pointer == 125 && y_pointer == 42)
||(x_pointer == 126 && y_pointer == 42)
||(x_pointer == 127 && y_pointer == 42)
||(x_pointer == 128 && y_pointer == 42)
||(x_pointer == 129 && y_pointer == 42)
||(x_pointer == 130 && y_pointer == 42)
||(x_pointer == 131 && y_pointer == 42)
||(x_pointer == 132 && y_pointer == 42)
||(x_pointer == 133 && y_pointer == 42)
||(x_pointer == 134 && y_pointer == 42)
||(x_pointer == 135 && y_pointer == 42)
||(x_pointer == 136 && y_pointer == 42)
||(x_pointer == 137 && y_pointer == 42)
||(x_pointer == 138 && y_pointer == 42)
||(x_pointer == 139 && y_pointer == 42)
||(x_pointer == 140 && y_pointer == 42)
||(x_pointer == 141 && y_pointer == 42)
||(x_pointer == 142 && y_pointer == 42)
||(x_pointer == 143 && y_pointer == 42)
||(x_pointer == 144 && y_pointer == 42)
||(x_pointer == 145 && y_pointer == 42)
||(x_pointer == 14 && y_pointer == 43)
||(x_pointer == 15 && y_pointer == 43)
||(x_pointer == 16 && y_pointer == 43)
||(x_pointer == 26 && y_pointer == 43)
||(x_pointer == 27 && y_pointer == 43)
||(x_pointer == 28 && y_pointer == 43)
||(x_pointer == 95 && y_pointer == 43)
||(x_pointer == 96 && y_pointer == 43)
||(x_pointer == 97 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 99 && y_pointer == 43)
||(x_pointer == 100 && y_pointer == 43)
||(x_pointer == 101 && y_pointer == 43)
||(x_pointer == 102 && y_pointer == 43)
||(x_pointer == 103 && y_pointer == 43)
||(x_pointer == 104 && y_pointer == 43)
||(x_pointer == 105 && y_pointer == 43)
||(x_pointer == 106 && y_pointer == 43)
||(x_pointer == 107 && y_pointer == 43)
||(x_pointer == 108 && y_pointer == 43)
||(x_pointer == 109 && y_pointer == 43)
||(x_pointer == 110 && y_pointer == 43)
||(x_pointer == 111 && y_pointer == 43)
||(x_pointer == 112 && y_pointer == 43)
||(x_pointer == 113 && y_pointer == 43)
||(x_pointer == 114 && y_pointer == 43)
||(x_pointer == 115 && y_pointer == 43)
||(x_pointer == 116 && y_pointer == 43)
||(x_pointer == 117 && y_pointer == 43)
||(x_pointer == 118 && y_pointer == 43)
||(x_pointer == 119 && y_pointer == 43)
||(x_pointer == 120 && y_pointer == 43)
||(x_pointer == 121 && y_pointer == 43)
||(x_pointer == 122 && y_pointer == 43)
||(x_pointer == 123 && y_pointer == 43)
||(x_pointer == 124 && y_pointer == 43)
||(x_pointer == 125 && y_pointer == 43)
||(x_pointer == 126 && y_pointer == 43)
||(x_pointer == 127 && y_pointer == 43)
||(x_pointer == 128 && y_pointer == 43)
||(x_pointer == 129 && y_pointer == 43)
||(x_pointer == 130 && y_pointer == 43)
||(x_pointer == 131 && y_pointer == 43)
||(x_pointer == 132 && y_pointer == 43)
||(x_pointer == 133 && y_pointer == 43)
||(x_pointer == 134 && y_pointer == 43)
||(x_pointer == 135 && y_pointer == 43)
||(x_pointer == 136 && y_pointer == 43)
||(x_pointer == 137 && y_pointer == 43)
||(x_pointer == 138 && y_pointer == 43)
||(x_pointer == 139 && y_pointer == 43)
||(x_pointer == 140 && y_pointer == 43)
||(x_pointer == 141 && y_pointer == 43)
||(x_pointer == 142 && y_pointer == 43)
||(x_pointer == 143 && y_pointer == 43)
||(x_pointer == 144 && y_pointer == 43)
||(x_pointer == 145 && y_pointer == 43)
||(x_pointer == 14 && y_pointer == 44)
||(x_pointer == 15 && y_pointer == 44)
||(x_pointer == 16 && y_pointer == 44)
||(x_pointer == 26 && y_pointer == 44)
||(x_pointer == 27 && y_pointer == 44)
||(x_pointer == 28 && y_pointer == 44)
||(x_pointer == 143 && y_pointer == 44)
||(x_pointer == 144 && y_pointer == 44)
||(x_pointer == 145 && y_pointer == 44)
||(x_pointer == 14 && y_pointer == 45)
||(x_pointer == 15 && y_pointer == 45)
||(x_pointer == 16 && y_pointer == 45)
||(x_pointer == 26 && y_pointer == 45)
||(x_pointer == 27 && y_pointer == 45)
||(x_pointer == 28 && y_pointer == 45)
||(x_pointer == 143 && y_pointer == 45)
||(x_pointer == 144 && y_pointer == 45)
||(x_pointer == 145 && y_pointer == 45)
||(x_pointer == 14 && y_pointer == 46)
||(x_pointer == 15 && y_pointer == 46)
||(x_pointer == 16 && y_pointer == 46)
||(x_pointer == 26 && y_pointer == 46)
||(x_pointer == 27 && y_pointer == 46)
||(x_pointer == 28 && y_pointer == 46)
||(x_pointer == 143 && y_pointer == 46)
||(x_pointer == 144 && y_pointer == 46)
||(x_pointer == 145 && y_pointer == 46)
||(x_pointer == 14 && y_pointer == 47)
||(x_pointer == 15 && y_pointer == 47)
||(x_pointer == 16 && y_pointer == 47)
||(x_pointer == 26 && y_pointer == 47)
||(x_pointer == 27 && y_pointer == 47)
||(x_pointer == 28 && y_pointer == 47)
||(x_pointer == 143 && y_pointer == 47)
||(x_pointer == 144 && y_pointer == 47)
||(x_pointer == 145 && y_pointer == 47)
||(x_pointer == 14 && y_pointer == 48)
||(x_pointer == 15 && y_pointer == 48)
||(x_pointer == 16 && y_pointer == 48)
||(x_pointer == 26 && y_pointer == 48)
||(x_pointer == 27 && y_pointer == 48)
||(x_pointer == 28 && y_pointer == 48)
||(x_pointer == 143 && y_pointer == 48)
||(x_pointer == 144 && y_pointer == 48)
||(x_pointer == 145 && y_pointer == 48)
||(x_pointer == 14 && y_pointer == 49)
||(x_pointer == 15 && y_pointer == 49)
||(x_pointer == 16 && y_pointer == 49)
||(x_pointer == 26 && y_pointer == 49)
||(x_pointer == 27 && y_pointer == 49)
||(x_pointer == 28 && y_pointer == 49)
||(x_pointer == 143 && y_pointer == 49)
||(x_pointer == 144 && y_pointer == 49)
||(x_pointer == 145 && y_pointer == 49)
||(x_pointer == 14 && y_pointer == 50)
||(x_pointer == 15 && y_pointer == 50)
||(x_pointer == 16 && y_pointer == 50)
||(x_pointer == 26 && y_pointer == 50)
||(x_pointer == 27 && y_pointer == 50)
||(x_pointer == 28 && y_pointer == 50)
||(x_pointer == 38 && y_pointer == 50)
||(x_pointer == 39 && y_pointer == 50)
||(x_pointer == 40 && y_pointer == 50)
||(x_pointer == 41 && y_pointer == 50)
||(x_pointer == 42 && y_pointer == 50)
||(x_pointer == 43 && y_pointer == 50)
||(x_pointer == 44 && y_pointer == 50)
||(x_pointer == 45 && y_pointer == 50)
||(x_pointer == 46 && y_pointer == 50)
||(x_pointer == 47 && y_pointer == 50)
||(x_pointer == 48 && y_pointer == 50)
||(x_pointer == 49 && y_pointer == 50)
||(x_pointer == 50 && y_pointer == 50)
||(x_pointer == 51 && y_pointer == 50)
||(x_pointer == 52 && y_pointer == 50)
||(x_pointer == 53 && y_pointer == 50)
||(x_pointer == 54 && y_pointer == 50)
||(x_pointer == 55 && y_pointer == 50)
||(x_pointer == 56 && y_pointer == 50)
||(x_pointer == 57 && y_pointer == 50)
||(x_pointer == 58 && y_pointer == 50)
||(x_pointer == 59 && y_pointer == 50)
||(x_pointer == 60 && y_pointer == 50)
||(x_pointer == 61 && y_pointer == 50)
||(x_pointer == 62 && y_pointer == 50)
||(x_pointer == 63 && y_pointer == 50)
||(x_pointer == 64 && y_pointer == 50)
||(x_pointer == 65 && y_pointer == 50)
||(x_pointer == 66 && y_pointer == 50)
||(x_pointer == 67 && y_pointer == 50)
||(x_pointer == 68 && y_pointer == 50)
||(x_pointer == 69 && y_pointer == 50)
||(x_pointer == 70 && y_pointer == 50)
||(x_pointer == 14 && y_pointer == 51)
||(x_pointer == 15 && y_pointer == 51)
||(x_pointer == 16 && y_pointer == 51)
||(x_pointer == 26 && y_pointer == 51)
||(x_pointer == 27 && y_pointer == 51)
||(x_pointer == 28 && y_pointer == 51)
||(x_pointer == 38 && y_pointer == 51)
||(x_pointer == 39 && y_pointer == 51)
||(x_pointer == 40 && y_pointer == 51)
||(x_pointer == 41 && y_pointer == 51)
||(x_pointer == 42 && y_pointer == 51)
||(x_pointer == 43 && y_pointer == 51)
||(x_pointer == 44 && y_pointer == 51)
||(x_pointer == 45 && y_pointer == 51)
||(x_pointer == 46 && y_pointer == 51)
||(x_pointer == 47 && y_pointer == 51)
||(x_pointer == 48 && y_pointer == 51)
||(x_pointer == 49 && y_pointer == 51)
||(x_pointer == 50 && y_pointer == 51)
||(x_pointer == 51 && y_pointer == 51)
||(x_pointer == 52 && y_pointer == 51)
||(x_pointer == 53 && y_pointer == 51)
||(x_pointer == 54 && y_pointer == 51)
||(x_pointer == 55 && y_pointer == 51)
||(x_pointer == 56 && y_pointer == 51)
||(x_pointer == 57 && y_pointer == 51)
||(x_pointer == 58 && y_pointer == 51)
||(x_pointer == 59 && y_pointer == 51)
||(x_pointer == 60 && y_pointer == 51)
||(x_pointer == 61 && y_pointer == 51)
||(x_pointer == 62 && y_pointer == 51)
||(x_pointer == 63 && y_pointer == 51)
||(x_pointer == 64 && y_pointer == 51)
||(x_pointer == 65 && y_pointer == 51)
||(x_pointer == 66 && y_pointer == 51)
||(x_pointer == 67 && y_pointer == 51)
||(x_pointer == 68 && y_pointer == 51)
||(x_pointer == 69 && y_pointer == 51)
||(x_pointer == 70 && y_pointer == 51)
||(x_pointer == 14 && y_pointer == 52)
||(x_pointer == 15 && y_pointer == 52)
||(x_pointer == 16 && y_pointer == 52)
||(x_pointer == 26 && y_pointer == 52)
||(x_pointer == 27 && y_pointer == 52)
||(x_pointer == 28 && y_pointer == 52)
||(x_pointer == 38 && y_pointer == 52)
||(x_pointer == 39 && y_pointer == 52)
||(x_pointer == 40 && y_pointer == 52)
||(x_pointer == 41 && y_pointer == 52)
||(x_pointer == 42 && y_pointer == 52)
||(x_pointer == 43 && y_pointer == 52)
||(x_pointer == 44 && y_pointer == 52)
||(x_pointer == 45 && y_pointer == 52)
||(x_pointer == 46 && y_pointer == 52)
||(x_pointer == 47 && y_pointer == 52)
||(x_pointer == 48 && y_pointer == 52)
||(x_pointer == 49 && y_pointer == 52)
||(x_pointer == 50 && y_pointer == 52)
||(x_pointer == 51 && y_pointer == 52)
||(x_pointer == 52 && y_pointer == 52)
||(x_pointer == 53 && y_pointer == 52)
||(x_pointer == 54 && y_pointer == 52)
||(x_pointer == 55 && y_pointer == 52)
||(x_pointer == 56 && y_pointer == 52)
||(x_pointer == 57 && y_pointer == 52)
||(x_pointer == 58 && y_pointer == 52)
||(x_pointer == 59 && y_pointer == 52)
||(x_pointer == 60 && y_pointer == 52)
||(x_pointer == 61 && y_pointer == 52)
||(x_pointer == 62 && y_pointer == 52)
||(x_pointer == 63 && y_pointer == 52)
||(x_pointer == 64 && y_pointer == 52)
||(x_pointer == 65 && y_pointer == 52)
||(x_pointer == 66 && y_pointer == 52)
||(x_pointer == 67 && y_pointer == 52)
||(x_pointer == 68 && y_pointer == 52)
||(x_pointer == 69 && y_pointer == 52)
||(x_pointer == 70 && y_pointer == 52)
||(x_pointer == 26 && y_pointer == 53)
||(x_pointer == 27 && y_pointer == 53)
||(x_pointer == 28 && y_pointer == 53)
||(x_pointer == 26 && y_pointer == 54)
||(x_pointer == 27 && y_pointer == 54)
||(x_pointer == 28 && y_pointer == 54)
||(x_pointer == 26 && y_pointer == 55)
||(x_pointer == 27 && y_pointer == 55)
||(x_pointer == 28 && y_pointer == 55)
||(x_pointer == 26 && y_pointer == 56)
||(x_pointer == 27 && y_pointer == 56)
||(x_pointer == 28 && y_pointer == 56)
||(x_pointer == 26 && y_pointer == 57)
||(x_pointer == 27 && y_pointer == 57)
||(x_pointer == 28 && y_pointer == 57)
||(x_pointer == 26 && y_pointer == 58)
||(x_pointer == 27 && y_pointer == 58)
||(x_pointer == 28 && y_pointer == 58)
||(x_pointer == 26 && y_pointer == 59)
||(x_pointer == 27 && y_pointer == 59)
||(x_pointer == 28 && y_pointer == 59)
||(x_pointer == 110 && y_pointer == 59)
||(x_pointer == 111 && y_pointer == 59)
||(x_pointer == 112 && y_pointer == 59)
||(x_pointer == 113 && y_pointer == 59)
||(x_pointer == 114 && y_pointer == 59)
||(x_pointer == 115 && y_pointer == 59)
||(x_pointer == 116 && y_pointer == 59)
||(x_pointer == 117 && y_pointer == 59)
||(x_pointer == 118 && y_pointer == 59)
||(x_pointer == 119 && y_pointer == 59)
||(x_pointer == 120 && y_pointer == 59)
||(x_pointer == 121 && y_pointer == 59)
||(x_pointer == 122 && y_pointer == 59)
||(x_pointer == 123 && y_pointer == 59)
||(x_pointer == 124 && y_pointer == 59)
||(x_pointer == 125 && y_pointer == 59)
||(x_pointer == 126 && y_pointer == 59)
||(x_pointer == 127 && y_pointer == 59)
||(x_pointer == 128 && y_pointer == 59)
||(x_pointer == 129 && y_pointer == 59)
||(x_pointer == 130 && y_pointer == 59)
||(x_pointer == 143 && y_pointer == 59)
||(x_pointer == 144 && y_pointer == 59)
||(x_pointer == 145 && y_pointer == 59)
||(x_pointer == 26 && y_pointer == 60)
||(x_pointer == 27 && y_pointer == 60)
||(x_pointer == 28 && y_pointer == 60)
||(x_pointer == 110 && y_pointer == 60)
||(x_pointer == 111 && y_pointer == 60)
||(x_pointer == 112 && y_pointer == 60)
||(x_pointer == 113 && y_pointer == 60)
||(x_pointer == 114 && y_pointer == 60)
||(x_pointer == 115 && y_pointer == 60)
||(x_pointer == 116 && y_pointer == 60)
||(x_pointer == 117 && y_pointer == 60)
||(x_pointer == 118 && y_pointer == 60)
||(x_pointer == 119 && y_pointer == 60)
||(x_pointer == 120 && y_pointer == 60)
||(x_pointer == 121 && y_pointer == 60)
||(x_pointer == 122 && y_pointer == 60)
||(x_pointer == 123 && y_pointer == 60)
||(x_pointer == 124 && y_pointer == 60)
||(x_pointer == 125 && y_pointer == 60)
||(x_pointer == 126 && y_pointer == 60)
||(x_pointer == 127 && y_pointer == 60)
||(x_pointer == 128 && y_pointer == 60)
||(x_pointer == 129 && y_pointer == 60)
||(x_pointer == 130 && y_pointer == 60)
||(x_pointer == 143 && y_pointer == 60)
||(x_pointer == 144 && y_pointer == 60)
||(x_pointer == 145 && y_pointer == 60)
||(x_pointer == 26 && y_pointer == 61)
||(x_pointer == 27 && y_pointer == 61)
||(x_pointer == 28 && y_pointer == 61)
||(x_pointer == 110 && y_pointer == 61)
||(x_pointer == 111 && y_pointer == 61)
||(x_pointer == 112 && y_pointer == 61)
||(x_pointer == 113 && y_pointer == 61)
||(x_pointer == 114 && y_pointer == 61)
||(x_pointer == 115 && y_pointer == 61)
||(x_pointer == 116 && y_pointer == 61)
||(x_pointer == 117 && y_pointer == 61)
||(x_pointer == 118 && y_pointer == 61)
||(x_pointer == 119 && y_pointer == 61)
||(x_pointer == 120 && y_pointer == 61)
||(x_pointer == 121 && y_pointer == 61)
||(x_pointer == 122 && y_pointer == 61)
||(x_pointer == 123 && y_pointer == 61)
||(x_pointer == 124 && y_pointer == 61)
||(x_pointer == 125 && y_pointer == 61)
||(x_pointer == 126 && y_pointer == 61)
||(x_pointer == 127 && y_pointer == 61)
||(x_pointer == 128 && y_pointer == 61)
||(x_pointer == 129 && y_pointer == 61)
||(x_pointer == 130 && y_pointer == 61)
||(x_pointer == 143 && y_pointer == 61)
||(x_pointer == 144 && y_pointer == 61)
||(x_pointer == 145 && y_pointer == 61)
||(x_pointer == 26 && y_pointer == 62)
||(x_pointer == 27 && y_pointer == 62)
||(x_pointer == 28 && y_pointer == 62)
||(x_pointer == 38 && y_pointer == 62)
||(x_pointer == 39 && y_pointer == 62)
||(x_pointer == 40 && y_pointer == 62)
||(x_pointer == 41 && y_pointer == 62)
||(x_pointer == 42 && y_pointer == 62)
||(x_pointer == 43 && y_pointer == 62)
||(x_pointer == 44 && y_pointer == 62)
||(x_pointer == 45 && y_pointer == 62)
||(x_pointer == 46 && y_pointer == 62)
||(x_pointer == 47 && y_pointer == 62)
||(x_pointer == 48 && y_pointer == 62)
||(x_pointer == 49 && y_pointer == 62)
||(x_pointer == 50 && y_pointer == 62)
||(x_pointer == 51 && y_pointer == 62)
||(x_pointer == 52 && y_pointer == 62)
||(x_pointer == 53 && y_pointer == 62)
||(x_pointer == 54 && y_pointer == 62)
||(x_pointer == 55 && y_pointer == 62)
||(x_pointer == 56 && y_pointer == 62)
||(x_pointer == 57 && y_pointer == 62)
||(x_pointer == 58 && y_pointer == 62)
||(x_pointer == 59 && y_pointer == 62)
||(x_pointer == 60 && y_pointer == 62)
||(x_pointer == 61 && y_pointer == 62)
||(x_pointer == 62 && y_pointer == 62)
||(x_pointer == 63 && y_pointer == 62)
||(x_pointer == 64 && y_pointer == 62)
||(x_pointer == 65 && y_pointer == 62)
||(x_pointer == 66 && y_pointer == 62)
||(x_pointer == 67 && y_pointer == 62)
||(x_pointer == 68 && y_pointer == 62)
||(x_pointer == 69 && y_pointer == 62)
||(x_pointer == 70 && y_pointer == 62)
||(x_pointer == 110 && y_pointer == 62)
||(x_pointer == 111 && y_pointer == 62)
||(x_pointer == 112 && y_pointer == 62)
||(x_pointer == 128 && y_pointer == 62)
||(x_pointer == 129 && y_pointer == 62)
||(x_pointer == 130 && y_pointer == 62)
||(x_pointer == 143 && y_pointer == 62)
||(x_pointer == 144 && y_pointer == 62)
||(x_pointer == 145 && y_pointer == 62)
||(x_pointer == 26 && y_pointer == 63)
||(x_pointer == 27 && y_pointer == 63)
||(x_pointer == 28 && y_pointer == 63)
||(x_pointer == 38 && y_pointer == 63)
||(x_pointer == 39 && y_pointer == 63)
||(x_pointer == 40 && y_pointer == 63)
||(x_pointer == 41 && y_pointer == 63)
||(x_pointer == 42 && y_pointer == 63)
||(x_pointer == 43 && y_pointer == 63)
||(x_pointer == 44 && y_pointer == 63)
||(x_pointer == 45 && y_pointer == 63)
||(x_pointer == 46 && y_pointer == 63)
||(x_pointer == 47 && y_pointer == 63)
||(x_pointer == 48 && y_pointer == 63)
||(x_pointer == 49 && y_pointer == 63)
||(x_pointer == 50 && y_pointer == 63)
||(x_pointer == 51 && y_pointer == 63)
||(x_pointer == 52 && y_pointer == 63)
||(x_pointer == 53 && y_pointer == 63)
||(x_pointer == 54 && y_pointer == 63)
||(x_pointer == 55 && y_pointer == 63)
||(x_pointer == 56 && y_pointer == 63)
||(x_pointer == 57 && y_pointer == 63)
||(x_pointer == 58 && y_pointer == 63)
||(x_pointer == 59 && y_pointer == 63)
||(x_pointer == 60 && y_pointer == 63)
||(x_pointer == 61 && y_pointer == 63)
||(x_pointer == 62 && y_pointer == 63)
||(x_pointer == 63 && y_pointer == 63)
||(x_pointer == 64 && y_pointer == 63)
||(x_pointer == 65 && y_pointer == 63)
||(x_pointer == 66 && y_pointer == 63)
||(x_pointer == 67 && y_pointer == 63)
||(x_pointer == 68 && y_pointer == 63)
||(x_pointer == 69 && y_pointer == 63)
||(x_pointer == 70 && y_pointer == 63)
||(x_pointer == 110 && y_pointer == 63)
||(x_pointer == 111 && y_pointer == 63)
||(x_pointer == 112 && y_pointer == 63)
||(x_pointer == 128 && y_pointer == 63)
||(x_pointer == 129 && y_pointer == 63)
||(x_pointer == 130 && y_pointer == 63)
||(x_pointer == 143 && y_pointer == 63)
||(x_pointer == 144 && y_pointer == 63)
||(x_pointer == 145 && y_pointer == 63)
||(x_pointer == 26 && y_pointer == 64)
||(x_pointer == 27 && y_pointer == 64)
||(x_pointer == 28 && y_pointer == 64)
||(x_pointer == 38 && y_pointer == 64)
||(x_pointer == 39 && y_pointer == 64)
||(x_pointer == 40 && y_pointer == 64)
||(x_pointer == 41 && y_pointer == 64)
||(x_pointer == 42 && y_pointer == 64)
||(x_pointer == 43 && y_pointer == 64)
||(x_pointer == 44 && y_pointer == 64)
||(x_pointer == 45 && y_pointer == 64)
||(x_pointer == 46 && y_pointer == 64)
||(x_pointer == 47 && y_pointer == 64)
||(x_pointer == 48 && y_pointer == 64)
||(x_pointer == 49 && y_pointer == 64)
||(x_pointer == 50 && y_pointer == 64)
||(x_pointer == 51 && y_pointer == 64)
||(x_pointer == 52 && y_pointer == 64)
||(x_pointer == 53 && y_pointer == 64)
||(x_pointer == 54 && y_pointer == 64)
||(x_pointer == 55 && y_pointer == 64)
||(x_pointer == 56 && y_pointer == 64)
||(x_pointer == 57 && y_pointer == 64)
||(x_pointer == 58 && y_pointer == 64)
||(x_pointer == 59 && y_pointer == 64)
||(x_pointer == 60 && y_pointer == 64)
||(x_pointer == 61 && y_pointer == 64)
||(x_pointer == 62 && y_pointer == 64)
||(x_pointer == 63 && y_pointer == 64)
||(x_pointer == 64 && y_pointer == 64)
||(x_pointer == 65 && y_pointer == 64)
||(x_pointer == 66 && y_pointer == 64)
||(x_pointer == 67 && y_pointer == 64)
||(x_pointer == 68 && y_pointer == 64)
||(x_pointer == 69 && y_pointer == 64)
||(x_pointer == 70 && y_pointer == 64)
||(x_pointer == 110 && y_pointer == 64)
||(x_pointer == 111 && y_pointer == 64)
||(x_pointer == 112 && y_pointer == 64)
||(x_pointer == 128 && y_pointer == 64)
||(x_pointer == 129 && y_pointer == 64)
||(x_pointer == 130 && y_pointer == 64)
||(x_pointer == 143 && y_pointer == 64)
||(x_pointer == 144 && y_pointer == 64)
||(x_pointer == 145 && y_pointer == 64)
||(x_pointer == 14 && y_pointer == 65)
||(x_pointer == 15 && y_pointer == 65)
||(x_pointer == 16 && y_pointer == 65)
||(x_pointer == 26 && y_pointer == 65)
||(x_pointer == 27 && y_pointer == 65)
||(x_pointer == 28 && y_pointer == 65)
||(x_pointer == 110 && y_pointer == 65)
||(x_pointer == 111 && y_pointer == 65)
||(x_pointer == 112 && y_pointer == 65)
||(x_pointer == 128 && y_pointer == 65)
||(x_pointer == 129 && y_pointer == 65)
||(x_pointer == 130 && y_pointer == 65)
||(x_pointer == 143 && y_pointer == 65)
||(x_pointer == 144 && y_pointer == 65)
||(x_pointer == 145 && y_pointer == 65)
||(x_pointer == 14 && y_pointer == 66)
||(x_pointer == 15 && y_pointer == 66)
||(x_pointer == 16 && y_pointer == 66)
||(x_pointer == 26 && y_pointer == 66)
||(x_pointer == 27 && y_pointer == 66)
||(x_pointer == 28 && y_pointer == 66)
||(x_pointer == 110 && y_pointer == 66)
||(x_pointer == 111 && y_pointer == 66)
||(x_pointer == 112 && y_pointer == 66)
||(x_pointer == 128 && y_pointer == 66)
||(x_pointer == 129 && y_pointer == 66)
||(x_pointer == 130 && y_pointer == 66)
||(x_pointer == 143 && y_pointer == 66)
||(x_pointer == 144 && y_pointer == 66)
||(x_pointer == 145 && y_pointer == 66)
||(x_pointer == 14 && y_pointer == 67)
||(x_pointer == 15 && y_pointer == 67)
||(x_pointer == 16 && y_pointer == 67)
||(x_pointer == 26 && y_pointer == 67)
||(x_pointer == 27 && y_pointer == 67)
||(x_pointer == 28 && y_pointer == 67)
||(x_pointer == 110 && y_pointer == 67)
||(x_pointer == 111 && y_pointer == 67)
||(x_pointer == 112 && y_pointer == 67)
||(x_pointer == 128 && y_pointer == 67)
||(x_pointer == 129 && y_pointer == 67)
||(x_pointer == 130 && y_pointer == 67)
||(x_pointer == 143 && y_pointer == 67)
||(x_pointer == 144 && y_pointer == 67)
||(x_pointer == 145 && y_pointer == 67)
||(x_pointer == 14 && y_pointer == 68)
||(x_pointer == 15 && y_pointer == 68)
||(x_pointer == 16 && y_pointer == 68)
||(x_pointer == 26 && y_pointer == 68)
||(x_pointer == 27 && y_pointer == 68)
||(x_pointer == 28 && y_pointer == 68)
||(x_pointer == 110 && y_pointer == 68)
||(x_pointer == 111 && y_pointer == 68)
||(x_pointer == 112 && y_pointer == 68)
||(x_pointer == 128 && y_pointer == 68)
||(x_pointer == 129 && y_pointer == 68)
||(x_pointer == 130 && y_pointer == 68)
||(x_pointer == 143 && y_pointer == 68)
||(x_pointer == 144 && y_pointer == 68)
||(x_pointer == 145 && y_pointer == 68)
||(x_pointer == 14 && y_pointer == 69)
||(x_pointer == 15 && y_pointer == 69)
||(x_pointer == 16 && y_pointer == 69)
||(x_pointer == 26 && y_pointer == 69)
||(x_pointer == 27 && y_pointer == 69)
||(x_pointer == 28 && y_pointer == 69)
||(x_pointer == 110 && y_pointer == 69)
||(x_pointer == 111 && y_pointer == 69)
||(x_pointer == 112 && y_pointer == 69)
||(x_pointer == 128 && y_pointer == 69)
||(x_pointer == 129 && y_pointer == 69)
||(x_pointer == 130 && y_pointer == 69)
||(x_pointer == 143 && y_pointer == 69)
||(x_pointer == 144 && y_pointer == 69)
||(x_pointer == 145 && y_pointer == 69)
||(x_pointer == 14 && y_pointer == 70)
||(x_pointer == 15 && y_pointer == 70)
||(x_pointer == 16 && y_pointer == 70)
||(x_pointer == 26 && y_pointer == 70)
||(x_pointer == 27 && y_pointer == 70)
||(x_pointer == 28 && y_pointer == 70)
||(x_pointer == 110 && y_pointer == 70)
||(x_pointer == 111 && y_pointer == 70)
||(x_pointer == 112 && y_pointer == 70)
||(x_pointer == 128 && y_pointer == 70)
||(x_pointer == 129 && y_pointer == 70)
||(x_pointer == 130 && y_pointer == 70)
||(x_pointer == 143 && y_pointer == 70)
||(x_pointer == 144 && y_pointer == 70)
||(x_pointer == 145 && y_pointer == 70)
||(x_pointer == 14 && y_pointer == 71)
||(x_pointer == 15 && y_pointer == 71)
||(x_pointer == 16 && y_pointer == 71)
||(x_pointer == 26 && y_pointer == 71)
||(x_pointer == 27 && y_pointer == 71)
||(x_pointer == 28 && y_pointer == 71)
||(x_pointer == 95 && y_pointer == 71)
||(x_pointer == 96 && y_pointer == 71)
||(x_pointer == 97 && y_pointer == 71)
||(x_pointer == 110 && y_pointer == 71)
||(x_pointer == 111 && y_pointer == 71)
||(x_pointer == 112 && y_pointer == 71)
||(x_pointer == 143 && y_pointer == 71)
||(x_pointer == 144 && y_pointer == 71)
||(x_pointer == 145 && y_pointer == 71)
||(x_pointer == 14 && y_pointer == 72)
||(x_pointer == 15 && y_pointer == 72)
||(x_pointer == 16 && y_pointer == 72)
||(x_pointer == 26 && y_pointer == 72)
||(x_pointer == 27 && y_pointer == 72)
||(x_pointer == 28 && y_pointer == 72)
||(x_pointer == 95 && y_pointer == 72)
||(x_pointer == 96 && y_pointer == 72)
||(x_pointer == 97 && y_pointer == 72)
||(x_pointer == 110 && y_pointer == 72)
||(x_pointer == 111 && y_pointer == 72)
||(x_pointer == 112 && y_pointer == 72)
||(x_pointer == 143 && y_pointer == 72)
||(x_pointer == 144 && y_pointer == 72)
||(x_pointer == 145 && y_pointer == 72)
||(x_pointer == 14 && y_pointer == 73)
||(x_pointer == 15 && y_pointer == 73)
||(x_pointer == 16 && y_pointer == 73)
||(x_pointer == 26 && y_pointer == 73)
||(x_pointer == 27 && y_pointer == 73)
||(x_pointer == 28 && y_pointer == 73)
||(x_pointer == 95 && y_pointer == 73)
||(x_pointer == 96 && y_pointer == 73)
||(x_pointer == 97 && y_pointer == 73)
||(x_pointer == 110 && y_pointer == 73)
||(x_pointer == 111 && y_pointer == 73)
||(x_pointer == 112 && y_pointer == 73)
||(x_pointer == 143 && y_pointer == 73)
||(x_pointer == 144 && y_pointer == 73)
||(x_pointer == 145 && y_pointer == 73)
||(x_pointer == 14 && y_pointer == 74)
||(x_pointer == 15 && y_pointer == 74)
||(x_pointer == 16 && y_pointer == 74)
||(x_pointer == 26 && y_pointer == 74)
||(x_pointer == 27 && y_pointer == 74)
||(x_pointer == 28 && y_pointer == 74)
||(x_pointer == 56 && y_pointer == 74)
||(x_pointer == 57 && y_pointer == 74)
||(x_pointer == 58 && y_pointer == 74)
||(x_pointer == 59 && y_pointer == 74)
||(x_pointer == 60 && y_pointer == 74)
||(x_pointer == 61 && y_pointer == 74)
||(x_pointer == 62 && y_pointer == 74)
||(x_pointer == 63 && y_pointer == 74)
||(x_pointer == 64 && y_pointer == 74)
||(x_pointer == 65 && y_pointer == 74)
||(x_pointer == 66 && y_pointer == 74)
||(x_pointer == 67 && y_pointer == 74)
||(x_pointer == 68 && y_pointer == 74)
||(x_pointer == 69 && y_pointer == 74)
||(x_pointer == 70 && y_pointer == 74)
||(x_pointer == 71 && y_pointer == 74)
||(x_pointer == 72 && y_pointer == 74)
||(x_pointer == 73 && y_pointer == 74)
||(x_pointer == 74 && y_pointer == 74)
||(x_pointer == 75 && y_pointer == 74)
||(x_pointer == 76 && y_pointer == 74)
||(x_pointer == 77 && y_pointer == 74)
||(x_pointer == 78 && y_pointer == 74)
||(x_pointer == 79 && y_pointer == 74)
||(x_pointer == 80 && y_pointer == 74)
||(x_pointer == 81 && y_pointer == 74)
||(x_pointer == 82 && y_pointer == 74)
||(x_pointer == 95 && y_pointer == 74)
||(x_pointer == 96 && y_pointer == 74)
||(x_pointer == 97 && y_pointer == 74)
||(x_pointer == 110 && y_pointer == 74)
||(x_pointer == 111 && y_pointer == 74)
||(x_pointer == 112 && y_pointer == 74)
||(x_pointer == 143 && y_pointer == 74)
||(x_pointer == 144 && y_pointer == 74)
||(x_pointer == 145 && y_pointer == 74)
||(x_pointer == 14 && y_pointer == 75)
||(x_pointer == 15 && y_pointer == 75)
||(x_pointer == 16 && y_pointer == 75)
||(x_pointer == 26 && y_pointer == 75)
||(x_pointer == 27 && y_pointer == 75)
||(x_pointer == 28 && y_pointer == 75)
||(x_pointer == 56 && y_pointer == 75)
||(x_pointer == 57 && y_pointer == 75)
||(x_pointer == 58 && y_pointer == 75)
||(x_pointer == 59 && y_pointer == 75)
||(x_pointer == 60 && y_pointer == 75)
||(x_pointer == 61 && y_pointer == 75)
||(x_pointer == 62 && y_pointer == 75)
||(x_pointer == 63 && y_pointer == 75)
||(x_pointer == 64 && y_pointer == 75)
||(x_pointer == 65 && y_pointer == 75)
||(x_pointer == 66 && y_pointer == 75)
||(x_pointer == 67 && y_pointer == 75)
||(x_pointer == 68 && y_pointer == 75)
||(x_pointer == 69 && y_pointer == 75)
||(x_pointer == 70 && y_pointer == 75)
||(x_pointer == 71 && y_pointer == 75)
||(x_pointer == 72 && y_pointer == 75)
||(x_pointer == 73 && y_pointer == 75)
||(x_pointer == 74 && y_pointer == 75)
||(x_pointer == 75 && y_pointer == 75)
||(x_pointer == 76 && y_pointer == 75)
||(x_pointer == 77 && y_pointer == 75)
||(x_pointer == 78 && y_pointer == 75)
||(x_pointer == 79 && y_pointer == 75)
||(x_pointer == 80 && y_pointer == 75)
||(x_pointer == 81 && y_pointer == 75)
||(x_pointer == 82 && y_pointer == 75)
||(x_pointer == 95 && y_pointer == 75)
||(x_pointer == 96 && y_pointer == 75)
||(x_pointer == 97 && y_pointer == 75)
||(x_pointer == 110 && y_pointer == 75)
||(x_pointer == 111 && y_pointer == 75)
||(x_pointer == 112 && y_pointer == 75)
||(x_pointer == 143 && y_pointer == 75)
||(x_pointer == 144 && y_pointer == 75)
||(x_pointer == 145 && y_pointer == 75)
||(x_pointer == 14 && y_pointer == 76)
||(x_pointer == 15 && y_pointer == 76)
||(x_pointer == 16 && y_pointer == 76)
||(x_pointer == 26 && y_pointer == 76)
||(x_pointer == 27 && y_pointer == 76)
||(x_pointer == 28 && y_pointer == 76)
||(x_pointer == 56 && y_pointer == 76)
||(x_pointer == 57 && y_pointer == 76)
||(x_pointer == 58 && y_pointer == 76)
||(x_pointer == 59 && y_pointer == 76)
||(x_pointer == 60 && y_pointer == 76)
||(x_pointer == 61 && y_pointer == 76)
||(x_pointer == 62 && y_pointer == 76)
||(x_pointer == 63 && y_pointer == 76)
||(x_pointer == 64 && y_pointer == 76)
||(x_pointer == 65 && y_pointer == 76)
||(x_pointer == 66 && y_pointer == 76)
||(x_pointer == 67 && y_pointer == 76)
||(x_pointer == 68 && y_pointer == 76)
||(x_pointer == 69 && y_pointer == 76)
||(x_pointer == 70 && y_pointer == 76)
||(x_pointer == 71 && y_pointer == 76)
||(x_pointer == 72 && y_pointer == 76)
||(x_pointer == 73 && y_pointer == 76)
||(x_pointer == 74 && y_pointer == 76)
||(x_pointer == 75 && y_pointer == 76)
||(x_pointer == 76 && y_pointer == 76)
||(x_pointer == 77 && y_pointer == 76)
||(x_pointer == 78 && y_pointer == 76)
||(x_pointer == 79 && y_pointer == 76)
||(x_pointer == 80 && y_pointer == 76)
||(x_pointer == 81 && y_pointer == 76)
||(x_pointer == 82 && y_pointer == 76)
||(x_pointer == 95 && y_pointer == 76)
||(x_pointer == 96 && y_pointer == 76)
||(x_pointer == 97 && y_pointer == 76)
||(x_pointer == 110 && y_pointer == 76)
||(x_pointer == 111 && y_pointer == 76)
||(x_pointer == 112 && y_pointer == 76)
||(x_pointer == 143 && y_pointer == 76)
||(x_pointer == 144 && y_pointer == 76)
||(x_pointer == 145 && y_pointer == 76)
||(x_pointer == 14 && y_pointer == 77)
||(x_pointer == 15 && y_pointer == 77)
||(x_pointer == 16 && y_pointer == 77)
||(x_pointer == 38 && y_pointer == 77)
||(x_pointer == 39 && y_pointer == 77)
||(x_pointer == 40 && y_pointer == 77)
||(x_pointer == 95 && y_pointer == 77)
||(x_pointer == 96 && y_pointer == 77)
||(x_pointer == 97 && y_pointer == 77)
||(x_pointer == 143 && y_pointer == 77)
||(x_pointer == 144 && y_pointer == 77)
||(x_pointer == 145 && y_pointer == 77)
||(x_pointer == 14 && y_pointer == 78)
||(x_pointer == 15 && y_pointer == 78)
||(x_pointer == 16 && y_pointer == 78)
||(x_pointer == 38 && y_pointer == 78)
||(x_pointer == 39 && y_pointer == 78)
||(x_pointer == 40 && y_pointer == 78)
||(x_pointer == 95 && y_pointer == 78)
||(x_pointer == 96 && y_pointer == 78)
||(x_pointer == 97 && y_pointer == 78)
||(x_pointer == 143 && y_pointer == 78)
||(x_pointer == 144 && y_pointer == 78)
||(x_pointer == 145 && y_pointer == 78)
||(x_pointer == 14 && y_pointer == 79)
||(x_pointer == 15 && y_pointer == 79)
||(x_pointer == 16 && y_pointer == 79)
||(x_pointer == 38 && y_pointer == 79)
||(x_pointer == 39 && y_pointer == 79)
||(x_pointer == 40 && y_pointer == 79)
||(x_pointer == 95 && y_pointer == 79)
||(x_pointer == 96 && y_pointer == 79)
||(x_pointer == 97 && y_pointer == 79)
||(x_pointer == 143 && y_pointer == 79)
||(x_pointer == 144 && y_pointer == 79)
||(x_pointer == 145 && y_pointer == 79)
||(x_pointer == 14 && y_pointer == 80)
||(x_pointer == 15 && y_pointer == 80)
||(x_pointer == 16 && y_pointer == 80)
||(x_pointer == 38 && y_pointer == 80)
||(x_pointer == 39 && y_pointer == 80)
||(x_pointer == 40 && y_pointer == 80)
||(x_pointer == 95 && y_pointer == 80)
||(x_pointer == 96 && y_pointer == 80)
||(x_pointer == 97 && y_pointer == 80)
||(x_pointer == 143 && y_pointer == 80)
||(x_pointer == 144 && y_pointer == 80)
||(x_pointer == 145 && y_pointer == 80)
||(x_pointer == 14 && y_pointer == 81)
||(x_pointer == 15 && y_pointer == 81)
||(x_pointer == 16 && y_pointer == 81)
||(x_pointer == 38 && y_pointer == 81)
||(x_pointer == 39 && y_pointer == 81)
||(x_pointer == 40 && y_pointer == 81)
||(x_pointer == 95 && y_pointer == 81)
||(x_pointer == 96 && y_pointer == 81)
||(x_pointer == 97 && y_pointer == 81)
||(x_pointer == 143 && y_pointer == 81)
||(x_pointer == 144 && y_pointer == 81)
||(x_pointer == 145 && y_pointer == 81)
||(x_pointer == 14 && y_pointer == 82)
||(x_pointer == 15 && y_pointer == 82)
||(x_pointer == 16 && y_pointer == 82)
||(x_pointer == 38 && y_pointer == 82)
||(x_pointer == 39 && y_pointer == 82)
||(x_pointer == 40 && y_pointer == 82)
||(x_pointer == 95 && y_pointer == 82)
||(x_pointer == 96 && y_pointer == 82)
||(x_pointer == 97 && y_pointer == 82)
||(x_pointer == 143 && y_pointer == 82)
||(x_pointer == 144 && y_pointer == 82)
||(x_pointer == 145 && y_pointer == 82)
||(x_pointer == 14 && y_pointer == 83)
||(x_pointer == 15 && y_pointer == 83)
||(x_pointer == 16 && y_pointer == 83)
||(x_pointer == 38 && y_pointer == 83)
||(x_pointer == 39 && y_pointer == 83)
||(x_pointer == 40 && y_pointer == 83)
||(x_pointer == 95 && y_pointer == 83)
||(x_pointer == 96 && y_pointer == 83)
||(x_pointer == 97 && y_pointer == 83)
||(x_pointer == 143 && y_pointer == 83)
||(x_pointer == 144 && y_pointer == 83)
||(x_pointer == 145 && y_pointer == 83)
||(x_pointer == 14 && y_pointer == 84)
||(x_pointer == 15 && y_pointer == 84)
||(x_pointer == 16 && y_pointer == 84)
||(x_pointer == 38 && y_pointer == 84)
||(x_pointer == 39 && y_pointer == 84)
||(x_pointer == 40 && y_pointer == 84)
||(x_pointer == 95 && y_pointer == 84)
||(x_pointer == 96 && y_pointer == 84)
||(x_pointer == 97 && y_pointer == 84)
||(x_pointer == 143 && y_pointer == 84)
||(x_pointer == 144 && y_pointer == 84)
||(x_pointer == 145 && y_pointer == 84)
||(x_pointer == 14 && y_pointer == 85)
||(x_pointer == 15 && y_pointer == 85)
||(x_pointer == 16 && y_pointer == 85)
||(x_pointer == 38 && y_pointer == 85)
||(x_pointer == 39 && y_pointer == 85)
||(x_pointer == 40 && y_pointer == 85)
||(x_pointer == 95 && y_pointer == 85)
||(x_pointer == 96 && y_pointer == 85)
||(x_pointer == 97 && y_pointer == 85)
||(x_pointer == 143 && y_pointer == 85)
||(x_pointer == 144 && y_pointer == 85)
||(x_pointer == 145 && y_pointer == 85)
||(x_pointer == 14 && y_pointer == 86)
||(x_pointer == 15 && y_pointer == 86)
||(x_pointer == 16 && y_pointer == 86)
||(x_pointer == 38 && y_pointer == 86)
||(x_pointer == 39 && y_pointer == 86)
||(x_pointer == 40 && y_pointer == 86)
||(x_pointer == 95 && y_pointer == 86)
||(x_pointer == 96 && y_pointer == 86)
||(x_pointer == 97 && y_pointer == 86)
||(x_pointer == 143 && y_pointer == 86)
||(x_pointer == 144 && y_pointer == 86)
||(x_pointer == 145 && y_pointer == 86)
||(x_pointer == 14 && y_pointer == 87)
||(x_pointer == 15 && y_pointer == 87)
||(x_pointer == 16 && y_pointer == 87)
||(x_pointer == 38 && y_pointer == 87)
||(x_pointer == 39 && y_pointer == 87)
||(x_pointer == 40 && y_pointer == 87)
||(x_pointer == 95 && y_pointer == 87)
||(x_pointer == 96 && y_pointer == 87)
||(x_pointer == 97 && y_pointer == 87)
||(x_pointer == 143 && y_pointer == 87)
||(x_pointer == 144 && y_pointer == 87)
||(x_pointer == 145 && y_pointer == 87)
||(x_pointer == 14 && y_pointer == 88)
||(x_pointer == 15 && y_pointer == 88)
||(x_pointer == 16 && y_pointer == 88)
||(x_pointer == 38 && y_pointer == 88)
||(x_pointer == 39 && y_pointer == 88)
||(x_pointer == 40 && y_pointer == 88)
||(x_pointer == 95 && y_pointer == 88)
||(x_pointer == 96 && y_pointer == 88)
||(x_pointer == 97 && y_pointer == 88)
||(x_pointer == 143 && y_pointer == 88)
||(x_pointer == 144 && y_pointer == 88)
||(x_pointer == 145 && y_pointer == 88)
||(x_pointer == 14 && y_pointer == 89)
||(x_pointer == 15 && y_pointer == 89)
||(x_pointer == 16 && y_pointer == 89)
||(x_pointer == 26 && y_pointer == 89)
||(x_pointer == 27 && y_pointer == 89)
||(x_pointer == 28 && y_pointer == 89)
||(x_pointer == 38 && y_pointer == 89)
||(x_pointer == 39 && y_pointer == 89)
||(x_pointer == 40 && y_pointer == 89)
||(x_pointer == 56 && y_pointer == 89)
||(x_pointer == 57 && y_pointer == 89)
||(x_pointer == 58 && y_pointer == 89)
||(x_pointer == 71 && y_pointer == 89)
||(x_pointer == 72 && y_pointer == 89)
||(x_pointer == 73 && y_pointer == 89)
||(x_pointer == 95 && y_pointer == 89)
||(x_pointer == 96 && y_pointer == 89)
||(x_pointer == 97 && y_pointer == 89)
||(x_pointer == 110 && y_pointer == 89)
||(x_pointer == 111 && y_pointer == 89)
||(x_pointer == 112 && y_pointer == 89)
||(x_pointer == 143 && y_pointer == 89)
||(x_pointer == 144 && y_pointer == 89)
||(x_pointer == 145 && y_pointer == 89)
||(x_pointer == 14 && y_pointer == 90)
||(x_pointer == 15 && y_pointer == 90)
||(x_pointer == 16 && y_pointer == 90)
||(x_pointer == 26 && y_pointer == 90)
||(x_pointer == 27 && y_pointer == 90)
||(x_pointer == 28 && y_pointer == 90)
||(x_pointer == 38 && y_pointer == 90)
||(x_pointer == 39 && y_pointer == 90)
||(x_pointer == 40 && y_pointer == 90)
||(x_pointer == 56 && y_pointer == 90)
||(x_pointer == 57 && y_pointer == 90)
||(x_pointer == 58 && y_pointer == 90)
||(x_pointer == 71 && y_pointer == 90)
||(x_pointer == 72 && y_pointer == 90)
||(x_pointer == 73 && y_pointer == 90)
||(x_pointer == 95 && y_pointer == 90)
||(x_pointer == 96 && y_pointer == 90)
||(x_pointer == 97 && y_pointer == 90)
||(x_pointer == 110 && y_pointer == 90)
||(x_pointer == 111 && y_pointer == 90)
||(x_pointer == 112 && y_pointer == 90)
||(x_pointer == 143 && y_pointer == 90)
||(x_pointer == 144 && y_pointer == 90)
||(x_pointer == 145 && y_pointer == 90)
||(x_pointer == 14 && y_pointer == 91)
||(x_pointer == 15 && y_pointer == 91)
||(x_pointer == 16 && y_pointer == 91)
||(x_pointer == 26 && y_pointer == 91)
||(x_pointer == 27 && y_pointer == 91)
||(x_pointer == 28 && y_pointer == 91)
||(x_pointer == 38 && y_pointer == 91)
||(x_pointer == 39 && y_pointer == 91)
||(x_pointer == 40 && y_pointer == 91)
||(x_pointer == 56 && y_pointer == 91)
||(x_pointer == 57 && y_pointer == 91)
||(x_pointer == 58 && y_pointer == 91)
||(x_pointer == 71 && y_pointer == 91)
||(x_pointer == 72 && y_pointer == 91)
||(x_pointer == 73 && y_pointer == 91)
||(x_pointer == 95 && y_pointer == 91)
||(x_pointer == 96 && y_pointer == 91)
||(x_pointer == 97 && y_pointer == 91)
||(x_pointer == 110 && y_pointer == 91)
||(x_pointer == 111 && y_pointer == 91)
||(x_pointer == 112 && y_pointer == 91)
||(x_pointer == 143 && y_pointer == 91)
||(x_pointer == 144 && y_pointer == 91)
||(x_pointer == 145 && y_pointer == 91)
||(x_pointer == 14 && y_pointer == 92)
||(x_pointer == 15 && y_pointer == 92)
||(x_pointer == 16 && y_pointer == 92)
||(x_pointer == 26 && y_pointer == 92)
||(x_pointer == 27 && y_pointer == 92)
||(x_pointer == 28 && y_pointer == 92)
||(x_pointer == 38 && y_pointer == 92)
||(x_pointer == 39 && y_pointer == 92)
||(x_pointer == 40 && y_pointer == 92)
||(x_pointer == 56 && y_pointer == 92)
||(x_pointer == 57 && y_pointer == 92)
||(x_pointer == 58 && y_pointer == 92)
||(x_pointer == 71 && y_pointer == 92)
||(x_pointer == 72 && y_pointer == 92)
||(x_pointer == 73 && y_pointer == 92)
||(x_pointer == 95 && y_pointer == 92)
||(x_pointer == 96 && y_pointer == 92)
||(x_pointer == 97 && y_pointer == 92)
||(x_pointer == 110 && y_pointer == 92)
||(x_pointer == 111 && y_pointer == 92)
||(x_pointer == 112 && y_pointer == 92)
||(x_pointer == 143 && y_pointer == 92)
||(x_pointer == 144 && y_pointer == 92)
||(x_pointer == 145 && y_pointer == 92)
||(x_pointer == 14 && y_pointer == 93)
||(x_pointer == 15 && y_pointer == 93)
||(x_pointer == 16 && y_pointer == 93)
||(x_pointer == 26 && y_pointer == 93)
||(x_pointer == 27 && y_pointer == 93)
||(x_pointer == 28 && y_pointer == 93)
||(x_pointer == 38 && y_pointer == 93)
||(x_pointer == 39 && y_pointer == 93)
||(x_pointer == 40 && y_pointer == 93)
||(x_pointer == 56 && y_pointer == 93)
||(x_pointer == 57 && y_pointer == 93)
||(x_pointer == 58 && y_pointer == 93)
||(x_pointer == 71 && y_pointer == 93)
||(x_pointer == 72 && y_pointer == 93)
||(x_pointer == 73 && y_pointer == 93)
||(x_pointer == 95 && y_pointer == 93)
||(x_pointer == 96 && y_pointer == 93)
||(x_pointer == 97 && y_pointer == 93)
||(x_pointer == 110 && y_pointer == 93)
||(x_pointer == 111 && y_pointer == 93)
||(x_pointer == 112 && y_pointer == 93)
||(x_pointer == 143 && y_pointer == 93)
||(x_pointer == 144 && y_pointer == 93)
||(x_pointer == 145 && y_pointer == 93)
||(x_pointer == 14 && y_pointer == 94)
||(x_pointer == 15 && y_pointer == 94)
||(x_pointer == 16 && y_pointer == 94)
||(x_pointer == 26 && y_pointer == 94)
||(x_pointer == 27 && y_pointer == 94)
||(x_pointer == 28 && y_pointer == 94)
||(x_pointer == 38 && y_pointer == 94)
||(x_pointer == 39 && y_pointer == 94)
||(x_pointer == 40 && y_pointer == 94)
||(x_pointer == 56 && y_pointer == 94)
||(x_pointer == 57 && y_pointer == 94)
||(x_pointer == 58 && y_pointer == 94)
||(x_pointer == 71 && y_pointer == 94)
||(x_pointer == 72 && y_pointer == 94)
||(x_pointer == 73 && y_pointer == 94)
||(x_pointer == 95 && y_pointer == 94)
||(x_pointer == 96 && y_pointer == 94)
||(x_pointer == 97 && y_pointer == 94)
||(x_pointer == 110 && y_pointer == 94)
||(x_pointer == 111 && y_pointer == 94)
||(x_pointer == 112 && y_pointer == 94)
||(x_pointer == 143 && y_pointer == 94)
||(x_pointer == 144 && y_pointer == 94)
||(x_pointer == 145 && y_pointer == 94)
||(x_pointer == 14 && y_pointer == 95)
||(x_pointer == 15 && y_pointer == 95)
||(x_pointer == 16 && y_pointer == 95)
||(x_pointer == 26 && y_pointer == 95)
||(x_pointer == 27 && y_pointer == 95)
||(x_pointer == 28 && y_pointer == 95)
||(x_pointer == 38 && y_pointer == 95)
||(x_pointer == 39 && y_pointer == 95)
||(x_pointer == 40 && y_pointer == 95)
||(x_pointer == 56 && y_pointer == 95)
||(x_pointer == 57 && y_pointer == 95)
||(x_pointer == 58 && y_pointer == 95)
||(x_pointer == 71 && y_pointer == 95)
||(x_pointer == 72 && y_pointer == 95)
||(x_pointer == 73 && y_pointer == 95)
||(x_pointer == 95 && y_pointer == 95)
||(x_pointer == 96 && y_pointer == 95)
||(x_pointer == 97 && y_pointer == 95)
||(x_pointer == 110 && y_pointer == 95)
||(x_pointer == 111 && y_pointer == 95)
||(x_pointer == 112 && y_pointer == 95)
||(x_pointer == 143 && y_pointer == 95)
||(x_pointer == 144 && y_pointer == 95)
||(x_pointer == 145 && y_pointer == 95)
||(x_pointer == 14 && y_pointer == 96)
||(x_pointer == 15 && y_pointer == 96)
||(x_pointer == 16 && y_pointer == 96)
||(x_pointer == 26 && y_pointer == 96)
||(x_pointer == 27 && y_pointer == 96)
||(x_pointer == 28 && y_pointer == 96)
||(x_pointer == 38 && y_pointer == 96)
||(x_pointer == 39 && y_pointer == 96)
||(x_pointer == 40 && y_pointer == 96)
||(x_pointer == 56 && y_pointer == 96)
||(x_pointer == 57 && y_pointer == 96)
||(x_pointer == 58 && y_pointer == 96)
||(x_pointer == 71 && y_pointer == 96)
||(x_pointer == 72 && y_pointer == 96)
||(x_pointer == 73 && y_pointer == 96)
||(x_pointer == 95 && y_pointer == 96)
||(x_pointer == 96 && y_pointer == 96)
||(x_pointer == 97 && y_pointer == 96)
||(x_pointer == 110 && y_pointer == 96)
||(x_pointer == 111 && y_pointer == 96)
||(x_pointer == 112 && y_pointer == 96)
||(x_pointer == 143 && y_pointer == 96)
||(x_pointer == 144 && y_pointer == 96)
||(x_pointer == 145 && y_pointer == 96)
||(x_pointer == 14 && y_pointer == 97)
||(x_pointer == 15 && y_pointer == 97)
||(x_pointer == 16 && y_pointer == 97)
||(x_pointer == 26 && y_pointer == 97)
||(x_pointer == 27 && y_pointer == 97)
||(x_pointer == 28 && y_pointer == 97)
||(x_pointer == 38 && y_pointer == 97)
||(x_pointer == 39 && y_pointer == 97)
||(x_pointer == 40 && y_pointer == 97)
||(x_pointer == 56 && y_pointer == 97)
||(x_pointer == 57 && y_pointer == 97)
||(x_pointer == 58 && y_pointer == 97)
||(x_pointer == 71 && y_pointer == 97)
||(x_pointer == 72 && y_pointer == 97)
||(x_pointer == 73 && y_pointer == 97)
||(x_pointer == 95 && y_pointer == 97)
||(x_pointer == 96 && y_pointer == 97)
||(x_pointer == 97 && y_pointer == 97)
||(x_pointer == 110 && y_pointer == 97)
||(x_pointer == 111 && y_pointer == 97)
||(x_pointer == 112 && y_pointer == 97)
||(x_pointer == 143 && y_pointer == 97)
||(x_pointer == 144 && y_pointer == 97)
||(x_pointer == 145 && y_pointer == 97)
||(x_pointer == 14 && y_pointer == 98)
||(x_pointer == 15 && y_pointer == 98)
||(x_pointer == 16 && y_pointer == 98)
||(x_pointer == 17 && y_pointer == 98)
||(x_pointer == 18 && y_pointer == 98)
||(x_pointer == 19 && y_pointer == 98)
||(x_pointer == 20 && y_pointer == 98)
||(x_pointer == 21 && y_pointer == 98)
||(x_pointer == 22 && y_pointer == 98)
||(x_pointer == 23 && y_pointer == 98)
||(x_pointer == 24 && y_pointer == 98)
||(x_pointer == 25 && y_pointer == 98)
||(x_pointer == 26 && y_pointer == 98)
||(x_pointer == 27 && y_pointer == 98)
||(x_pointer == 28 && y_pointer == 98)
||(x_pointer == 38 && y_pointer == 98)
||(x_pointer == 39 && y_pointer == 98)
||(x_pointer == 40 && y_pointer == 98)
||(x_pointer == 41 && y_pointer == 98)
||(x_pointer == 42 && y_pointer == 98)
||(x_pointer == 43 && y_pointer == 98)
||(x_pointer == 44 && y_pointer == 98)
||(x_pointer == 45 && y_pointer == 98)
||(x_pointer == 46 && y_pointer == 98)
||(x_pointer == 47 && y_pointer == 98)
||(x_pointer == 48 && y_pointer == 98)
||(x_pointer == 49 && y_pointer == 98)
||(x_pointer == 50 && y_pointer == 98)
||(x_pointer == 51 && y_pointer == 98)
||(x_pointer == 52 && y_pointer == 98)
||(x_pointer == 53 && y_pointer == 98)
||(x_pointer == 54 && y_pointer == 98)
||(x_pointer == 55 && y_pointer == 98)
||(x_pointer == 56 && y_pointer == 98)
||(x_pointer == 57 && y_pointer == 98)
||(x_pointer == 58 && y_pointer == 98)
||(x_pointer == 71 && y_pointer == 98)
||(x_pointer == 72 && y_pointer == 98)
||(x_pointer == 73 && y_pointer == 98)
||(x_pointer == 74 && y_pointer == 98)
||(x_pointer == 75 && y_pointer == 98)
||(x_pointer == 76 && y_pointer == 98)
||(x_pointer == 77 && y_pointer == 98)
||(x_pointer == 78 && y_pointer == 98)
||(x_pointer == 79 && y_pointer == 98)
||(x_pointer == 80 && y_pointer == 98)
||(x_pointer == 81 && y_pointer == 98)
||(x_pointer == 82 && y_pointer == 98)
||(x_pointer == 83 && y_pointer == 98)
||(x_pointer == 84 && y_pointer == 98)
||(x_pointer == 85 && y_pointer == 98)
||(x_pointer == 86 && y_pointer == 98)
||(x_pointer == 87 && y_pointer == 98)
||(x_pointer == 88 && y_pointer == 98)
||(x_pointer == 89 && y_pointer == 98)
||(x_pointer == 90 && y_pointer == 98)
||(x_pointer == 91 && y_pointer == 98)
||(x_pointer == 92 && y_pointer == 98)
||(x_pointer == 93 && y_pointer == 98)
||(x_pointer == 94 && y_pointer == 98)
||(x_pointer == 95 && y_pointer == 98)
||(x_pointer == 96 && y_pointer == 98)
||(x_pointer == 97 && y_pointer == 98)
||(x_pointer == 110 && y_pointer == 98)
||(x_pointer == 111 && y_pointer == 98)
||(x_pointer == 112 && y_pointer == 98)
||(x_pointer == 113 && y_pointer == 98)
||(x_pointer == 114 && y_pointer == 98)
||(x_pointer == 115 && y_pointer == 98)
||(x_pointer == 116 && y_pointer == 98)
||(x_pointer == 117 && y_pointer == 98)
||(x_pointer == 118 && y_pointer == 98)
||(x_pointer == 119 && y_pointer == 98)
||(x_pointer == 120 && y_pointer == 98)
||(x_pointer == 121 && y_pointer == 98)
||(x_pointer == 122 && y_pointer == 98)
||(x_pointer == 123 && y_pointer == 98)
||(x_pointer == 124 && y_pointer == 98)
||(x_pointer == 125 && y_pointer == 98)
||(x_pointer == 126 && y_pointer == 98)
||(x_pointer == 127 && y_pointer == 98)
||(x_pointer == 128 && y_pointer == 98)
||(x_pointer == 129 && y_pointer == 98)
||(x_pointer == 130 && y_pointer == 98)
||(x_pointer == 131 && y_pointer == 98)
||(x_pointer == 132 && y_pointer == 98)
||(x_pointer == 133 && y_pointer == 98)
||(x_pointer == 134 && y_pointer == 98)
||(x_pointer == 135 && y_pointer == 98)
||(x_pointer == 136 && y_pointer == 98)
||(x_pointer == 137 && y_pointer == 98)
||(x_pointer == 138 && y_pointer == 98)
||(x_pointer == 139 && y_pointer == 98)
||(x_pointer == 140 && y_pointer == 98)
||(x_pointer == 141 && y_pointer == 98)
||(x_pointer == 142 && y_pointer == 98)
||(x_pointer == 143 && y_pointer == 98)
||(x_pointer == 144 && y_pointer == 98)
||(x_pointer == 145 && y_pointer == 98)
||(x_pointer == 14 && y_pointer == 99)
||(x_pointer == 15 && y_pointer == 99)
||(x_pointer == 16 && y_pointer == 99)
||(x_pointer == 17 && y_pointer == 99)
||(x_pointer == 18 && y_pointer == 99)
||(x_pointer == 19 && y_pointer == 99)
||(x_pointer == 20 && y_pointer == 99)
||(x_pointer == 21 && y_pointer == 99)
||(x_pointer == 22 && y_pointer == 99)
||(x_pointer == 23 && y_pointer == 99)
||(x_pointer == 24 && y_pointer == 99)
||(x_pointer == 25 && y_pointer == 99)
||(x_pointer == 26 && y_pointer == 99)
||(x_pointer == 27 && y_pointer == 99)
||(x_pointer == 28 && y_pointer == 99)
||(x_pointer == 38 && y_pointer == 99)
||(x_pointer == 39 && y_pointer == 99)
||(x_pointer == 40 && y_pointer == 99)
||(x_pointer == 41 && y_pointer == 99)
||(x_pointer == 42 && y_pointer == 99)
||(x_pointer == 43 && y_pointer == 99)
||(x_pointer == 44 && y_pointer == 99)
||(x_pointer == 45 && y_pointer == 99)
||(x_pointer == 46 && y_pointer == 99)
||(x_pointer == 47 && y_pointer == 99)
||(x_pointer == 48 && y_pointer == 99)
||(x_pointer == 49 && y_pointer == 99)
||(x_pointer == 50 && y_pointer == 99)
||(x_pointer == 51 && y_pointer == 99)
||(x_pointer == 52 && y_pointer == 99)
||(x_pointer == 53 && y_pointer == 99)
||(x_pointer == 54 && y_pointer == 99)
||(x_pointer == 55 && y_pointer == 99)
||(x_pointer == 56 && y_pointer == 99)
||(x_pointer == 57 && y_pointer == 99)
||(x_pointer == 58 && y_pointer == 99)
||(x_pointer == 71 && y_pointer == 99)
||(x_pointer == 72 && y_pointer == 99)
||(x_pointer == 73 && y_pointer == 99)
||(x_pointer == 74 && y_pointer == 99)
||(x_pointer == 75 && y_pointer == 99)
||(x_pointer == 76 && y_pointer == 99)
||(x_pointer == 77 && y_pointer == 99)
||(x_pointer == 78 && y_pointer == 99)
||(x_pointer == 79 && y_pointer == 99)
||(x_pointer == 80 && y_pointer == 99)
||(x_pointer == 81 && y_pointer == 99)
||(x_pointer == 82 && y_pointer == 99)
||(x_pointer == 83 && y_pointer == 99)
||(x_pointer == 84 && y_pointer == 99)
||(x_pointer == 85 && y_pointer == 99)
||(x_pointer == 86 && y_pointer == 99)
||(x_pointer == 87 && y_pointer == 99)
||(x_pointer == 88 && y_pointer == 99)
||(x_pointer == 89 && y_pointer == 99)
||(x_pointer == 90 && y_pointer == 99)
||(x_pointer == 91 && y_pointer == 99)
||(x_pointer == 92 && y_pointer == 99)
||(x_pointer == 93 && y_pointer == 99)
||(x_pointer == 94 && y_pointer == 99)
||(x_pointer == 95 && y_pointer == 99)
||(x_pointer == 96 && y_pointer == 99)
||(x_pointer == 97 && y_pointer == 99)
||(x_pointer == 110 && y_pointer == 99)
||(x_pointer == 111 && y_pointer == 99)
||(x_pointer == 112 && y_pointer == 99)
||(x_pointer == 113 && y_pointer == 99)
||(x_pointer == 114 && y_pointer == 99)
||(x_pointer == 115 && y_pointer == 99)
||(x_pointer == 116 && y_pointer == 99)
||(x_pointer == 117 && y_pointer == 99)
||(x_pointer == 118 && y_pointer == 99)
||(x_pointer == 119 && y_pointer == 99)
||(x_pointer == 120 && y_pointer == 99)
||(x_pointer == 121 && y_pointer == 99)
||(x_pointer == 122 && y_pointer == 99)
||(x_pointer == 123 && y_pointer == 99)
||(x_pointer == 124 && y_pointer == 99)
||(x_pointer == 125 && y_pointer == 99)
||(x_pointer == 126 && y_pointer == 99)
||(x_pointer == 127 && y_pointer == 99)
||(x_pointer == 128 && y_pointer == 99)
||(x_pointer == 129 && y_pointer == 99)
||(x_pointer == 130 && y_pointer == 99)
||(x_pointer == 131 && y_pointer == 99)
||(x_pointer == 132 && y_pointer == 99)
||(x_pointer == 133 && y_pointer == 99)
||(x_pointer == 134 && y_pointer == 99)
||(x_pointer == 135 && y_pointer == 99)
||(x_pointer == 136 && y_pointer == 99)
||(x_pointer == 137 && y_pointer == 99)
||(x_pointer == 138 && y_pointer == 99)
||(x_pointer == 139 && y_pointer == 99)
||(x_pointer == 140 && y_pointer == 99)
||(x_pointer == 141 && y_pointer == 99)
||(x_pointer == 142 && y_pointer == 99)
||(x_pointer == 143 && y_pointer == 99)
||(x_pointer == 144 && y_pointer == 99)
||(x_pointer == 145 && y_pointer == 99)
||(x_pointer == 14 && y_pointer == 100)
||(x_pointer == 15 && y_pointer == 100)
||(x_pointer == 16 && y_pointer == 100)
||(x_pointer == 17 && y_pointer == 100)
||(x_pointer == 18 && y_pointer == 100)
||(x_pointer == 19 && y_pointer == 100)
||(x_pointer == 20 && y_pointer == 100)
||(x_pointer == 21 && y_pointer == 100)
||(x_pointer == 22 && y_pointer == 100)
||(x_pointer == 23 && y_pointer == 100)
||(x_pointer == 24 && y_pointer == 100)
||(x_pointer == 25 && y_pointer == 100)
||(x_pointer == 26 && y_pointer == 100)
||(x_pointer == 27 && y_pointer == 100)
||(x_pointer == 28 && y_pointer == 100)
||(x_pointer == 38 && y_pointer == 100)
||(x_pointer == 39 && y_pointer == 100)
||(x_pointer == 40 && y_pointer == 100)
||(x_pointer == 41 && y_pointer == 100)
||(x_pointer == 42 && y_pointer == 100)
||(x_pointer == 43 && y_pointer == 100)
||(x_pointer == 44 && y_pointer == 100)
||(x_pointer == 45 && y_pointer == 100)
||(x_pointer == 46 && y_pointer == 100)
||(x_pointer == 47 && y_pointer == 100)
||(x_pointer == 48 && y_pointer == 100)
||(x_pointer == 49 && y_pointer == 100)
||(x_pointer == 50 && y_pointer == 100)
||(x_pointer == 51 && y_pointer == 100)
||(x_pointer == 52 && y_pointer == 100)
||(x_pointer == 53 && y_pointer == 100)
||(x_pointer == 54 && y_pointer == 100)
||(x_pointer == 55 && y_pointer == 100)
||(x_pointer == 56 && y_pointer == 100)
||(x_pointer == 57 && y_pointer == 100)
||(x_pointer == 58 && y_pointer == 100)
||(x_pointer == 71 && y_pointer == 100)
||(x_pointer == 72 && y_pointer == 100)
||(x_pointer == 73 && y_pointer == 100)
||(x_pointer == 74 && y_pointer == 100)
||(x_pointer == 75 && y_pointer == 100)
||(x_pointer == 76 && y_pointer == 100)
||(x_pointer == 77 && y_pointer == 100)
||(x_pointer == 78 && y_pointer == 100)
||(x_pointer == 79 && y_pointer == 100)
||(x_pointer == 80 && y_pointer == 100)
||(x_pointer == 81 && y_pointer == 100)
||(x_pointer == 82 && y_pointer == 100)
||(x_pointer == 83 && y_pointer == 100)
||(x_pointer == 84 && y_pointer == 100)
||(x_pointer == 85 && y_pointer == 100)
||(x_pointer == 86 && y_pointer == 100)
||(x_pointer == 87 && y_pointer == 100)
||(x_pointer == 88 && y_pointer == 100)
||(x_pointer == 89 && y_pointer == 100)
||(x_pointer == 90 && y_pointer == 100)
||(x_pointer == 91 && y_pointer == 100)
||(x_pointer == 92 && y_pointer == 100)
||(x_pointer == 93 && y_pointer == 100)
||(x_pointer == 94 && y_pointer == 100)
||(x_pointer == 95 && y_pointer == 100)
||(x_pointer == 96 && y_pointer == 100)
||(x_pointer == 97 && y_pointer == 100)
||(x_pointer == 110 && y_pointer == 100)
||(x_pointer == 111 && y_pointer == 100)
||(x_pointer == 112 && y_pointer == 100)
||(x_pointer == 113 && y_pointer == 100)
||(x_pointer == 114 && y_pointer == 100)
||(x_pointer == 115 && y_pointer == 100)
||(x_pointer == 116 && y_pointer == 100)
||(x_pointer == 117 && y_pointer == 100)
||(x_pointer == 118 && y_pointer == 100)
||(x_pointer == 119 && y_pointer == 100)
||(x_pointer == 120 && y_pointer == 100)
||(x_pointer == 121 && y_pointer == 100)
||(x_pointer == 122 && y_pointer == 100)
||(x_pointer == 123 && y_pointer == 100)
||(x_pointer == 124 && y_pointer == 100)
||(x_pointer == 125 && y_pointer == 100)
||(x_pointer == 126 && y_pointer == 100)
||(x_pointer == 127 && y_pointer == 100)
||(x_pointer == 128 && y_pointer == 100)
||(x_pointer == 129 && y_pointer == 100)
||(x_pointer == 130 && y_pointer == 100)
||(x_pointer == 131 && y_pointer == 100)
||(x_pointer == 132 && y_pointer == 100)
||(x_pointer == 133 && y_pointer == 100)
||(x_pointer == 134 && y_pointer == 100)
||(x_pointer == 135 && y_pointer == 100)
||(x_pointer == 136 && y_pointer == 100)
||(x_pointer == 137 && y_pointer == 100)
||(x_pointer == 138 && y_pointer == 100)
||(x_pointer == 139 && y_pointer == 100)
||(x_pointer == 140 && y_pointer == 100)
||(x_pointer == 141 && y_pointer == 100)
||(x_pointer == 142 && y_pointer == 100)
||(x_pointer == 143 && y_pointer == 100)
||(x_pointer == 144 && y_pointer == 100)
||(x_pointer == 145 && y_pointer == 100));
	
	wire barrier_pixel_7 = current_level == 7 && ((x_pointer == 36 && y_pointer == 23)
||(x_pointer == 37 && y_pointer == 23)
||(x_pointer == 38 && y_pointer == 23)
||(x_pointer == 39 && y_pointer == 23)
||(x_pointer == 40 && y_pointer == 23)
||(x_pointer == 41 && y_pointer == 23)
||(x_pointer == 42 && y_pointer == 23)
||(x_pointer == 43 && y_pointer == 23)
||(x_pointer == 44 && y_pointer == 23)
||(x_pointer == 45 && y_pointer == 23)
||(x_pointer == 46 && y_pointer == 23)
||(x_pointer == 47 && y_pointer == 23)
||(x_pointer == 48 && y_pointer == 23)
||(x_pointer == 49 && y_pointer == 23)
||(x_pointer == 50 && y_pointer == 23)
||(x_pointer == 51 && y_pointer == 23)
||(x_pointer == 52 && y_pointer == 23)
||(x_pointer == 53 && y_pointer == 23)
||(x_pointer == 54 && y_pointer == 23)
||(x_pointer == 55 && y_pointer == 23)
||(x_pointer == 56 && y_pointer == 23)
||(x_pointer == 57 && y_pointer == 23)
||(x_pointer == 58 && y_pointer == 23)
||(x_pointer == 59 && y_pointer == 23)
||(x_pointer == 60 && y_pointer == 23)
||(x_pointer == 67 && y_pointer == 23)
||(x_pointer == 68 && y_pointer == 23)
||(x_pointer == 69 && y_pointer == 23)
||(x_pointer == 70 && y_pointer == 23)
||(x_pointer == 71 && y_pointer == 23)
||(x_pointer == 72 && y_pointer == 23)
||(x_pointer == 73 && y_pointer == 23)
||(x_pointer == 74 && y_pointer == 23)
||(x_pointer == 75 && y_pointer == 23)
||(x_pointer == 76 && y_pointer == 23)
||(x_pointer == 77 && y_pointer == 23)
||(x_pointer == 78 && y_pointer == 23)
||(x_pointer == 79 && y_pointer == 23)
||(x_pointer == 80 && y_pointer == 23)
||(x_pointer == 81 && y_pointer == 23)
||(x_pointer == 82 && y_pointer == 23)
||(x_pointer == 83 && y_pointer == 23)
||(x_pointer == 84 && y_pointer == 23)
||(x_pointer == 85 && y_pointer == 23)
||(x_pointer == 86 && y_pointer == 23)
||(x_pointer == 87 && y_pointer == 23)
||(x_pointer == 88 && y_pointer == 23)
||(x_pointer == 89 && y_pointer == 23)
||(x_pointer == 96 && y_pointer == 23)
||(x_pointer == 97 && y_pointer == 23)
||(x_pointer == 98 && y_pointer == 23)
||(x_pointer == 99 && y_pointer == 23)
||(x_pointer == 100 && y_pointer == 23)
||(x_pointer == 101 && y_pointer == 23)
||(x_pointer == 102 && y_pointer == 23)
||(x_pointer == 103 && y_pointer == 23)
||(x_pointer == 104 && y_pointer == 23)
||(x_pointer == 105 && y_pointer == 23)
||(x_pointer == 106 && y_pointer == 23)
||(x_pointer == 107 && y_pointer == 23)
||(x_pointer == 108 && y_pointer == 23)
||(x_pointer == 109 && y_pointer == 23)
||(x_pointer == 110 && y_pointer == 23)
||(x_pointer == 111 && y_pointer == 23)
||(x_pointer == 112 && y_pointer == 23)
||(x_pointer == 113 && y_pointer == 23)
||(x_pointer == 114 && y_pointer == 23)
||(x_pointer == 115 && y_pointer == 23)
||(x_pointer == 116 && y_pointer == 23)
||(x_pointer == 117 && y_pointer == 23)
||(x_pointer == 118 && y_pointer == 23)
||(x_pointer == 119 && y_pointer == 23)
||(x_pointer == 120 && y_pointer == 23)
||(x_pointer == 36 && y_pointer == 24)
||(x_pointer == 37 && y_pointer == 24)
||(x_pointer == 38 && y_pointer == 24)
||(x_pointer == 39 && y_pointer == 24)
||(x_pointer == 40 && y_pointer == 24)
||(x_pointer == 41 && y_pointer == 24)
||(x_pointer == 42 && y_pointer == 24)
||(x_pointer == 43 && y_pointer == 24)
||(x_pointer == 44 && y_pointer == 24)
||(x_pointer == 45 && y_pointer == 24)
||(x_pointer == 46 && y_pointer == 24)
||(x_pointer == 47 && y_pointer == 24)
||(x_pointer == 48 && y_pointer == 24)
||(x_pointer == 49 && y_pointer == 24)
||(x_pointer == 50 && y_pointer == 24)
||(x_pointer == 51 && y_pointer == 24)
||(x_pointer == 52 && y_pointer == 24)
||(x_pointer == 53 && y_pointer == 24)
||(x_pointer == 54 && y_pointer == 24)
||(x_pointer == 55 && y_pointer == 24)
||(x_pointer == 56 && y_pointer == 24)
||(x_pointer == 57 && y_pointer == 24)
||(x_pointer == 58 && y_pointer == 24)
||(x_pointer == 59 && y_pointer == 24)
||(x_pointer == 60 && y_pointer == 24)
||(x_pointer == 67 && y_pointer == 24)
||(x_pointer == 68 && y_pointer == 24)
||(x_pointer == 69 && y_pointer == 24)
||(x_pointer == 70 && y_pointer == 24)
||(x_pointer == 71 && y_pointer == 24)
||(x_pointer == 72 && y_pointer == 24)
||(x_pointer == 73 && y_pointer == 24)
||(x_pointer == 74 && y_pointer == 24)
||(x_pointer == 75 && y_pointer == 24)
||(x_pointer == 76 && y_pointer == 24)
||(x_pointer == 77 && y_pointer == 24)
||(x_pointer == 78 && y_pointer == 24)
||(x_pointer == 79 && y_pointer == 24)
||(x_pointer == 80 && y_pointer == 24)
||(x_pointer == 81 && y_pointer == 24)
||(x_pointer == 82 && y_pointer == 24)
||(x_pointer == 83 && y_pointer == 24)
||(x_pointer == 84 && y_pointer == 24)
||(x_pointer == 85 && y_pointer == 24)
||(x_pointer == 86 && y_pointer == 24)
||(x_pointer == 87 && y_pointer == 24)
||(x_pointer == 88 && y_pointer == 24)
||(x_pointer == 89 && y_pointer == 24)
||(x_pointer == 96 && y_pointer == 24)
||(x_pointer == 97 && y_pointer == 24)
||(x_pointer == 98 && y_pointer == 24)
||(x_pointer == 99 && y_pointer == 24)
||(x_pointer == 100 && y_pointer == 24)
||(x_pointer == 101 && y_pointer == 24)
||(x_pointer == 102 && y_pointer == 24)
||(x_pointer == 103 && y_pointer == 24)
||(x_pointer == 104 && y_pointer == 24)
||(x_pointer == 105 && y_pointer == 24)
||(x_pointer == 106 && y_pointer == 24)
||(x_pointer == 107 && y_pointer == 24)
||(x_pointer == 108 && y_pointer == 24)
||(x_pointer == 109 && y_pointer == 24)
||(x_pointer == 110 && y_pointer == 24)
||(x_pointer == 111 && y_pointer == 24)
||(x_pointer == 112 && y_pointer == 24)
||(x_pointer == 113 && y_pointer == 24)
||(x_pointer == 114 && y_pointer == 24)
||(x_pointer == 115 && y_pointer == 24)
||(x_pointer == 116 && y_pointer == 24)
||(x_pointer == 117 && y_pointer == 24)
||(x_pointer == 118 && y_pointer == 24)
||(x_pointer == 119 && y_pointer == 24)
||(x_pointer == 120 && y_pointer == 24)
||(x_pointer == 36 && y_pointer == 25)
||(x_pointer == 37 && y_pointer == 25)
||(x_pointer == 38 && y_pointer == 25)
||(x_pointer == 39 && y_pointer == 25)
||(x_pointer == 40 && y_pointer == 25)
||(x_pointer == 41 && y_pointer == 25)
||(x_pointer == 42 && y_pointer == 25)
||(x_pointer == 43 && y_pointer == 25)
||(x_pointer == 44 && y_pointer == 25)
||(x_pointer == 45 && y_pointer == 25)
||(x_pointer == 46 && y_pointer == 25)
||(x_pointer == 47 && y_pointer == 25)
||(x_pointer == 48 && y_pointer == 25)
||(x_pointer == 49 && y_pointer == 25)
||(x_pointer == 50 && y_pointer == 25)
||(x_pointer == 51 && y_pointer == 25)
||(x_pointer == 52 && y_pointer == 25)
||(x_pointer == 53 && y_pointer == 25)
||(x_pointer == 54 && y_pointer == 25)
||(x_pointer == 55 && y_pointer == 25)
||(x_pointer == 56 && y_pointer == 25)
||(x_pointer == 57 && y_pointer == 25)
||(x_pointer == 58 && y_pointer == 25)
||(x_pointer == 59 && y_pointer == 25)
||(x_pointer == 60 && y_pointer == 25)
||(x_pointer == 67 && y_pointer == 25)
||(x_pointer == 68 && y_pointer == 25)
||(x_pointer == 69 && y_pointer == 25)
||(x_pointer == 70 && y_pointer == 25)
||(x_pointer == 71 && y_pointer == 25)
||(x_pointer == 72 && y_pointer == 25)
||(x_pointer == 73 && y_pointer == 25)
||(x_pointer == 74 && y_pointer == 25)
||(x_pointer == 75 && y_pointer == 25)
||(x_pointer == 76 && y_pointer == 25)
||(x_pointer == 77 && y_pointer == 25)
||(x_pointer == 78 && y_pointer == 25)
||(x_pointer == 79 && y_pointer == 25)
||(x_pointer == 80 && y_pointer == 25)
||(x_pointer == 81 && y_pointer == 25)
||(x_pointer == 82 && y_pointer == 25)
||(x_pointer == 83 && y_pointer == 25)
||(x_pointer == 84 && y_pointer == 25)
||(x_pointer == 85 && y_pointer == 25)
||(x_pointer == 86 && y_pointer == 25)
||(x_pointer == 87 && y_pointer == 25)
||(x_pointer == 88 && y_pointer == 25)
||(x_pointer == 89 && y_pointer == 25)
||(x_pointer == 96 && y_pointer == 25)
||(x_pointer == 97 && y_pointer == 25)
||(x_pointer == 98 && y_pointer == 25)
||(x_pointer == 99 && y_pointer == 25)
||(x_pointer == 100 && y_pointer == 25)
||(x_pointer == 101 && y_pointer == 25)
||(x_pointer == 102 && y_pointer == 25)
||(x_pointer == 103 && y_pointer == 25)
||(x_pointer == 104 && y_pointer == 25)
||(x_pointer == 105 && y_pointer == 25)
||(x_pointer == 106 && y_pointer == 25)
||(x_pointer == 107 && y_pointer == 25)
||(x_pointer == 108 && y_pointer == 25)
||(x_pointer == 109 && y_pointer == 25)
||(x_pointer == 110 && y_pointer == 25)
||(x_pointer == 111 && y_pointer == 25)
||(x_pointer == 112 && y_pointer == 25)
||(x_pointer == 113 && y_pointer == 25)
||(x_pointer == 114 && y_pointer == 25)
||(x_pointer == 115 && y_pointer == 25)
||(x_pointer == 116 && y_pointer == 25)
||(x_pointer == 117 && y_pointer == 25)
||(x_pointer == 118 && y_pointer == 25)
||(x_pointer == 119 && y_pointer == 25)
||(x_pointer == 120 && y_pointer == 25)
||(x_pointer == 36 && y_pointer == 26)
||(x_pointer == 37 && y_pointer == 26)
||(x_pointer == 38 && y_pointer == 26)
||(x_pointer == 39 && y_pointer == 26)
||(x_pointer == 40 && y_pointer == 26)
||(x_pointer == 41 && y_pointer == 26)
||(x_pointer == 42 && y_pointer == 26)
||(x_pointer == 43 && y_pointer == 26)
||(x_pointer == 44 && y_pointer == 26)
||(x_pointer == 45 && y_pointer == 26)
||(x_pointer == 46 && y_pointer == 26)
||(x_pointer == 47 && y_pointer == 26)
||(x_pointer == 48 && y_pointer == 26)
||(x_pointer == 49 && y_pointer == 26)
||(x_pointer == 50 && y_pointer == 26)
||(x_pointer == 51 && y_pointer == 26)
||(x_pointer == 52 && y_pointer == 26)
||(x_pointer == 53 && y_pointer == 26)
||(x_pointer == 54 && y_pointer == 26)
||(x_pointer == 55 && y_pointer == 26)
||(x_pointer == 56 && y_pointer == 26)
||(x_pointer == 57 && y_pointer == 26)
||(x_pointer == 58 && y_pointer == 26)
||(x_pointer == 59 && y_pointer == 26)
||(x_pointer == 60 && y_pointer == 26)
||(x_pointer == 67 && y_pointer == 26)
||(x_pointer == 68 && y_pointer == 26)
||(x_pointer == 69 && y_pointer == 26)
||(x_pointer == 70 && y_pointer == 26)
||(x_pointer == 71 && y_pointer == 26)
||(x_pointer == 72 && y_pointer == 26)
||(x_pointer == 73 && y_pointer == 26)
||(x_pointer == 74 && y_pointer == 26)
||(x_pointer == 75 && y_pointer == 26)
||(x_pointer == 76 && y_pointer == 26)
||(x_pointer == 77 && y_pointer == 26)
||(x_pointer == 78 && y_pointer == 26)
||(x_pointer == 79 && y_pointer == 26)
||(x_pointer == 80 && y_pointer == 26)
||(x_pointer == 81 && y_pointer == 26)
||(x_pointer == 82 && y_pointer == 26)
||(x_pointer == 83 && y_pointer == 26)
||(x_pointer == 84 && y_pointer == 26)
||(x_pointer == 85 && y_pointer == 26)
||(x_pointer == 86 && y_pointer == 26)
||(x_pointer == 87 && y_pointer == 26)
||(x_pointer == 88 && y_pointer == 26)
||(x_pointer == 89 && y_pointer == 26)
||(x_pointer == 96 && y_pointer == 26)
||(x_pointer == 97 && y_pointer == 26)
||(x_pointer == 98 && y_pointer == 26)
||(x_pointer == 99 && y_pointer == 26)
||(x_pointer == 100 && y_pointer == 26)
||(x_pointer == 101 && y_pointer == 26)
||(x_pointer == 102 && y_pointer == 26)
||(x_pointer == 103 && y_pointer == 26)
||(x_pointer == 104 && y_pointer == 26)
||(x_pointer == 105 && y_pointer == 26)
||(x_pointer == 106 && y_pointer == 26)
||(x_pointer == 107 && y_pointer == 26)
||(x_pointer == 108 && y_pointer == 26)
||(x_pointer == 109 && y_pointer == 26)
||(x_pointer == 110 && y_pointer == 26)
||(x_pointer == 111 && y_pointer == 26)
||(x_pointer == 112 && y_pointer == 26)
||(x_pointer == 113 && y_pointer == 26)
||(x_pointer == 114 && y_pointer == 26)
||(x_pointer == 115 && y_pointer == 26)
||(x_pointer == 116 && y_pointer == 26)
||(x_pointer == 117 && y_pointer == 26)
||(x_pointer == 118 && y_pointer == 26)
||(x_pointer == 119 && y_pointer == 26)
||(x_pointer == 120 && y_pointer == 26)
||(x_pointer == 36 && y_pointer == 27)
||(x_pointer == 37 && y_pointer == 27)
||(x_pointer == 38 && y_pointer == 27)
||(x_pointer == 39 && y_pointer == 27)
||(x_pointer == 67 && y_pointer == 27)
||(x_pointer == 68 && y_pointer == 27)
||(x_pointer == 69 && y_pointer == 27)
||(x_pointer == 70 && y_pointer == 27)
||(x_pointer == 86 && y_pointer == 27)
||(x_pointer == 87 && y_pointer == 27)
||(x_pointer == 88 && y_pointer == 27)
||(x_pointer == 89 && y_pointer == 27)
||(x_pointer == 96 && y_pointer == 27)
||(x_pointer == 97 && y_pointer == 27)
||(x_pointer == 98 && y_pointer == 27)
||(x_pointer == 99 && y_pointer == 27)
||(x_pointer == 36 && y_pointer == 28)
||(x_pointer == 37 && y_pointer == 28)
||(x_pointer == 38 && y_pointer == 28)
||(x_pointer == 39 && y_pointer == 28)
||(x_pointer == 67 && y_pointer == 28)
||(x_pointer == 68 && y_pointer == 28)
||(x_pointer == 69 && y_pointer == 28)
||(x_pointer == 70 && y_pointer == 28)
||(x_pointer == 86 && y_pointer == 28)
||(x_pointer == 87 && y_pointer == 28)
||(x_pointer == 88 && y_pointer == 28)
||(x_pointer == 89 && y_pointer == 28)
||(x_pointer == 96 && y_pointer == 28)
||(x_pointer == 97 && y_pointer == 28)
||(x_pointer == 98 && y_pointer == 28)
||(x_pointer == 99 && y_pointer == 28)
||(x_pointer == 36 && y_pointer == 29)
||(x_pointer == 37 && y_pointer == 29)
||(x_pointer == 38 && y_pointer == 29)
||(x_pointer == 39 && y_pointer == 29)
||(x_pointer == 67 && y_pointer == 29)
||(x_pointer == 68 && y_pointer == 29)
||(x_pointer == 69 && y_pointer == 29)
||(x_pointer == 70 && y_pointer == 29)
||(x_pointer == 96 && y_pointer == 29)
||(x_pointer == 97 && y_pointer == 29)
||(x_pointer == 98 && y_pointer == 29)
||(x_pointer == 99 && y_pointer == 29)
||(x_pointer == 36 && y_pointer == 30)
||(x_pointer == 37 && y_pointer == 30)
||(x_pointer == 38 && y_pointer == 30)
||(x_pointer == 39 && y_pointer == 30)
||(x_pointer == 67 && y_pointer == 30)
||(x_pointer == 68 && y_pointer == 30)
||(x_pointer == 69 && y_pointer == 30)
||(x_pointer == 70 && y_pointer == 30)
||(x_pointer == 96 && y_pointer == 30)
||(x_pointer == 97 && y_pointer == 30)
||(x_pointer == 98 && y_pointer == 30)
||(x_pointer == 99 && y_pointer == 30)
||(x_pointer == 36 && y_pointer == 31)
||(x_pointer == 37 && y_pointer == 31)
||(x_pointer == 38 && y_pointer == 31)
||(x_pointer == 39 && y_pointer == 31)
||(x_pointer == 67 && y_pointer == 31)
||(x_pointer == 68 && y_pointer == 31)
||(x_pointer == 69 && y_pointer == 31)
||(x_pointer == 70 && y_pointer == 31)
||(x_pointer == 96 && y_pointer == 31)
||(x_pointer == 97 && y_pointer == 31)
||(x_pointer == 98 && y_pointer == 31)
||(x_pointer == 99 && y_pointer == 31)
||(x_pointer == 36 && y_pointer == 32)
||(x_pointer == 37 && y_pointer == 32)
||(x_pointer == 38 && y_pointer == 32)
||(x_pointer == 39 && y_pointer == 32)
||(x_pointer == 67 && y_pointer == 32)
||(x_pointer == 68 && y_pointer == 32)
||(x_pointer == 69 && y_pointer == 32)
||(x_pointer == 70 && y_pointer == 32)
||(x_pointer == 96 && y_pointer == 32)
||(x_pointer == 97 && y_pointer == 32)
||(x_pointer == 98 && y_pointer == 32)
||(x_pointer == 99 && y_pointer == 32)
||(x_pointer == 36 && y_pointer == 33)
||(x_pointer == 37 && y_pointer == 33)
||(x_pointer == 38 && y_pointer == 33)
||(x_pointer == 39 && y_pointer == 33)
||(x_pointer == 67 && y_pointer == 33)
||(x_pointer == 68 && y_pointer == 33)
||(x_pointer == 69 && y_pointer == 33)
||(x_pointer == 70 && y_pointer == 33)
||(x_pointer == 96 && y_pointer == 33)
||(x_pointer == 97 && y_pointer == 33)
||(x_pointer == 98 && y_pointer == 33)
||(x_pointer == 99 && y_pointer == 33)
||(x_pointer == 36 && y_pointer == 34)
||(x_pointer == 37 && y_pointer == 34)
||(x_pointer == 38 && y_pointer == 34)
||(x_pointer == 39 && y_pointer == 34)
||(x_pointer == 67 && y_pointer == 34)
||(x_pointer == 68 && y_pointer == 34)
||(x_pointer == 69 && y_pointer == 34)
||(x_pointer == 70 && y_pointer == 34)
||(x_pointer == 96 && y_pointer == 34)
||(x_pointer == 97 && y_pointer == 34)
||(x_pointer == 98 && y_pointer == 34)
||(x_pointer == 99 && y_pointer == 34)
||(x_pointer == 36 && y_pointer == 35)
||(x_pointer == 37 && y_pointer == 35)
||(x_pointer == 38 && y_pointer == 35)
||(x_pointer == 39 && y_pointer == 35)
||(x_pointer == 67 && y_pointer == 35)
||(x_pointer == 68 && y_pointer == 35)
||(x_pointer == 69 && y_pointer == 35)
||(x_pointer == 70 && y_pointer == 35)
||(x_pointer == 96 && y_pointer == 35)
||(x_pointer == 97 && y_pointer == 35)
||(x_pointer == 98 && y_pointer == 35)
||(x_pointer == 99 && y_pointer == 35)
||(x_pointer == 36 && y_pointer == 36)
||(x_pointer == 37 && y_pointer == 36)
||(x_pointer == 38 && y_pointer == 36)
||(x_pointer == 39 && y_pointer == 36)
||(x_pointer == 67 && y_pointer == 36)
||(x_pointer == 68 && y_pointer == 36)
||(x_pointer == 69 && y_pointer == 36)
||(x_pointer == 70 && y_pointer == 36)
||(x_pointer == 71 && y_pointer == 36)
||(x_pointer == 72 && y_pointer == 36)
||(x_pointer == 73 && y_pointer == 36)
||(x_pointer == 74 && y_pointer == 36)
||(x_pointer == 75 && y_pointer == 36)
||(x_pointer == 76 && y_pointer == 36)
||(x_pointer == 77 && y_pointer == 36)
||(x_pointer == 78 && y_pointer == 36)
||(x_pointer == 79 && y_pointer == 36)
||(x_pointer == 80 && y_pointer == 36)
||(x_pointer == 81 && y_pointer == 36)
||(x_pointer == 82 && y_pointer == 36)
||(x_pointer == 83 && y_pointer == 36)
||(x_pointer == 84 && y_pointer == 36)
||(x_pointer == 85 && y_pointer == 36)
||(x_pointer == 86 && y_pointer == 36)
||(x_pointer == 87 && y_pointer == 36)
||(x_pointer == 88 && y_pointer == 36)
||(x_pointer == 89 && y_pointer == 36)
||(x_pointer == 96 && y_pointer == 36)
||(x_pointer == 97 && y_pointer == 36)
||(x_pointer == 98 && y_pointer == 36)
||(x_pointer == 99 && y_pointer == 36)
||(x_pointer == 36 && y_pointer == 37)
||(x_pointer == 37 && y_pointer == 37)
||(x_pointer == 38 && y_pointer == 37)
||(x_pointer == 39 && y_pointer == 37)
||(x_pointer == 67 && y_pointer == 37)
||(x_pointer == 68 && y_pointer == 37)
||(x_pointer == 69 && y_pointer == 37)
||(x_pointer == 70 && y_pointer == 37)
||(x_pointer == 71 && y_pointer == 37)
||(x_pointer == 72 && y_pointer == 37)
||(x_pointer == 73 && y_pointer == 37)
||(x_pointer == 74 && y_pointer == 37)
||(x_pointer == 75 && y_pointer == 37)
||(x_pointer == 76 && y_pointer == 37)
||(x_pointer == 77 && y_pointer == 37)
||(x_pointer == 78 && y_pointer == 37)
||(x_pointer == 79 && y_pointer == 37)
||(x_pointer == 80 && y_pointer == 37)
||(x_pointer == 81 && y_pointer == 37)
||(x_pointer == 82 && y_pointer == 37)
||(x_pointer == 83 && y_pointer == 37)
||(x_pointer == 84 && y_pointer == 37)
||(x_pointer == 85 && y_pointer == 37)
||(x_pointer == 86 && y_pointer == 37)
||(x_pointer == 87 && y_pointer == 37)
||(x_pointer == 88 && y_pointer == 37)
||(x_pointer == 89 && y_pointer == 37)
||(x_pointer == 96 && y_pointer == 37)
||(x_pointer == 97 && y_pointer == 37)
||(x_pointer == 98 && y_pointer == 37)
||(x_pointer == 99 && y_pointer == 37)
||(x_pointer == 36 && y_pointer == 38)
||(x_pointer == 37 && y_pointer == 38)
||(x_pointer == 38 && y_pointer == 38)
||(x_pointer == 39 && y_pointer == 38)
||(x_pointer == 67 && y_pointer == 38)
||(x_pointer == 68 && y_pointer == 38)
||(x_pointer == 69 && y_pointer == 38)
||(x_pointer == 70 && y_pointer == 38)
||(x_pointer == 71 && y_pointer == 38)
||(x_pointer == 72 && y_pointer == 38)
||(x_pointer == 73 && y_pointer == 38)
||(x_pointer == 74 && y_pointer == 38)
||(x_pointer == 75 && y_pointer == 38)
||(x_pointer == 76 && y_pointer == 38)
||(x_pointer == 77 && y_pointer == 38)
||(x_pointer == 78 && y_pointer == 38)
||(x_pointer == 79 && y_pointer == 38)
||(x_pointer == 80 && y_pointer == 38)
||(x_pointer == 81 && y_pointer == 38)
||(x_pointer == 82 && y_pointer == 38)
||(x_pointer == 83 && y_pointer == 38)
||(x_pointer == 84 && y_pointer == 38)
||(x_pointer == 85 && y_pointer == 38)
||(x_pointer == 86 && y_pointer == 38)
||(x_pointer == 87 && y_pointer == 38)
||(x_pointer == 88 && y_pointer == 38)
||(x_pointer == 89 && y_pointer == 38)
||(x_pointer == 96 && y_pointer == 38)
||(x_pointer == 97 && y_pointer == 38)
||(x_pointer == 98 && y_pointer == 38)
||(x_pointer == 99 && y_pointer == 38)
||(x_pointer == 36 && y_pointer == 39)
||(x_pointer == 37 && y_pointer == 39)
||(x_pointer == 38 && y_pointer == 39)
||(x_pointer == 39 && y_pointer == 39)
||(x_pointer == 67 && y_pointer == 39)
||(x_pointer == 68 && y_pointer == 39)
||(x_pointer == 69 && y_pointer == 39)
||(x_pointer == 70 && y_pointer == 39)
||(x_pointer == 71 && y_pointer == 39)
||(x_pointer == 72 && y_pointer == 39)
||(x_pointer == 73 && y_pointer == 39)
||(x_pointer == 74 && y_pointer == 39)
||(x_pointer == 75 && y_pointer == 39)
||(x_pointer == 76 && y_pointer == 39)
||(x_pointer == 77 && y_pointer == 39)
||(x_pointer == 78 && y_pointer == 39)
||(x_pointer == 79 && y_pointer == 39)
||(x_pointer == 80 && y_pointer == 39)
||(x_pointer == 81 && y_pointer == 39)
||(x_pointer == 82 && y_pointer == 39)
||(x_pointer == 83 && y_pointer == 39)
||(x_pointer == 84 && y_pointer == 39)
||(x_pointer == 85 && y_pointer == 39)
||(x_pointer == 86 && y_pointer == 39)
||(x_pointer == 87 && y_pointer == 39)
||(x_pointer == 88 && y_pointer == 39)
||(x_pointer == 89 && y_pointer == 39)
||(x_pointer == 96 && y_pointer == 39)
||(x_pointer == 97 && y_pointer == 39)
||(x_pointer == 98 && y_pointer == 39)
||(x_pointer == 99 && y_pointer == 39)
||(x_pointer == 36 && y_pointer == 40)
||(x_pointer == 37 && y_pointer == 40)
||(x_pointer == 38 && y_pointer == 40)
||(x_pointer == 39 && y_pointer == 40)
||(x_pointer == 86 && y_pointer == 40)
||(x_pointer == 87 && y_pointer == 40)
||(x_pointer == 88 && y_pointer == 40)
||(x_pointer == 89 && y_pointer == 40)
||(x_pointer == 96 && y_pointer == 40)
||(x_pointer == 97 && y_pointer == 40)
||(x_pointer == 98 && y_pointer == 40)
||(x_pointer == 99 && y_pointer == 40)
||(x_pointer == 36 && y_pointer == 41)
||(x_pointer == 37 && y_pointer == 41)
||(x_pointer == 38 && y_pointer == 41)
||(x_pointer == 39 && y_pointer == 41)
||(x_pointer == 86 && y_pointer == 41)
||(x_pointer == 87 && y_pointer == 41)
||(x_pointer == 88 && y_pointer == 41)
||(x_pointer == 89 && y_pointer == 41)
||(x_pointer == 96 && y_pointer == 41)
||(x_pointer == 97 && y_pointer == 41)
||(x_pointer == 98 && y_pointer == 41)
||(x_pointer == 99 && y_pointer == 41)
||(x_pointer == 36 && y_pointer == 42)
||(x_pointer == 37 && y_pointer == 42)
||(x_pointer == 38 && y_pointer == 42)
||(x_pointer == 39 && y_pointer == 42)
||(x_pointer == 86 && y_pointer == 42)
||(x_pointer == 87 && y_pointer == 42)
||(x_pointer == 88 && y_pointer == 42)
||(x_pointer == 89 && y_pointer == 42)
||(x_pointer == 96 && y_pointer == 42)
||(x_pointer == 97 && y_pointer == 42)
||(x_pointer == 98 && y_pointer == 42)
||(x_pointer == 99 && y_pointer == 42)
||(x_pointer == 36 && y_pointer == 43)
||(x_pointer == 37 && y_pointer == 43)
||(x_pointer == 38 && y_pointer == 43)
||(x_pointer == 39 && y_pointer == 43)
||(x_pointer == 86 && y_pointer == 43)
||(x_pointer == 87 && y_pointer == 43)
||(x_pointer == 88 && y_pointer == 43)
||(x_pointer == 89 && y_pointer == 43)
||(x_pointer == 96 && y_pointer == 43)
||(x_pointer == 97 && y_pointer == 43)
||(x_pointer == 98 && y_pointer == 43)
||(x_pointer == 99 && y_pointer == 43)
||(x_pointer == 36 && y_pointer == 44)
||(x_pointer == 37 && y_pointer == 44)
||(x_pointer == 38 && y_pointer == 44)
||(x_pointer == 39 && y_pointer == 44)
||(x_pointer == 86 && y_pointer == 44)
||(x_pointer == 87 && y_pointer == 44)
||(x_pointer == 88 && y_pointer == 44)
||(x_pointer == 89 && y_pointer == 44)
||(x_pointer == 96 && y_pointer == 44)
||(x_pointer == 97 && y_pointer == 44)
||(x_pointer == 98 && y_pointer == 44)
||(x_pointer == 99 && y_pointer == 44)
||(x_pointer == 36 && y_pointer == 45)
||(x_pointer == 37 && y_pointer == 45)
||(x_pointer == 38 && y_pointer == 45)
||(x_pointer == 39 && y_pointer == 45)
||(x_pointer == 86 && y_pointer == 45)
||(x_pointer == 87 && y_pointer == 45)
||(x_pointer == 88 && y_pointer == 45)
||(x_pointer == 89 && y_pointer == 45)
||(x_pointer == 96 && y_pointer == 45)
||(x_pointer == 97 && y_pointer == 45)
||(x_pointer == 98 && y_pointer == 45)
||(x_pointer == 99 && y_pointer == 45)
||(x_pointer == 36 && y_pointer == 46)
||(x_pointer == 37 && y_pointer == 46)
||(x_pointer == 38 && y_pointer == 46)
||(x_pointer == 39 && y_pointer == 46)
||(x_pointer == 86 && y_pointer == 46)
||(x_pointer == 87 && y_pointer == 46)
||(x_pointer == 88 && y_pointer == 46)
||(x_pointer == 89 && y_pointer == 46)
||(x_pointer == 96 && y_pointer == 46)
||(x_pointer == 97 && y_pointer == 46)
||(x_pointer == 98 && y_pointer == 46)
||(x_pointer == 99 && y_pointer == 46)
||(x_pointer == 36 && y_pointer == 47)
||(x_pointer == 37 && y_pointer == 47)
||(x_pointer == 38 && y_pointer == 47)
||(x_pointer == 39 && y_pointer == 47)
||(x_pointer == 67 && y_pointer == 47)
||(x_pointer == 68 && y_pointer == 47)
||(x_pointer == 69 && y_pointer == 47)
||(x_pointer == 70 && y_pointer == 47)
||(x_pointer == 86 && y_pointer == 47)
||(x_pointer == 87 && y_pointer == 47)
||(x_pointer == 88 && y_pointer == 47)
||(x_pointer == 89 && y_pointer == 47)
||(x_pointer == 96 && y_pointer == 47)
||(x_pointer == 97 && y_pointer == 47)
||(x_pointer == 98 && y_pointer == 47)
||(x_pointer == 99 && y_pointer == 47)
||(x_pointer == 36 && y_pointer == 48)
||(x_pointer == 37 && y_pointer == 48)
||(x_pointer == 38 && y_pointer == 48)
||(x_pointer == 39 && y_pointer == 48)
||(x_pointer == 67 && y_pointer == 48)
||(x_pointer == 68 && y_pointer == 48)
||(x_pointer == 69 && y_pointer == 48)
||(x_pointer == 70 && y_pointer == 48)
||(x_pointer == 86 && y_pointer == 48)
||(x_pointer == 87 && y_pointer == 48)
||(x_pointer == 88 && y_pointer == 48)
||(x_pointer == 89 && y_pointer == 48)
||(x_pointer == 96 && y_pointer == 48)
||(x_pointer == 97 && y_pointer == 48)
||(x_pointer == 98 && y_pointer == 48)
||(x_pointer == 99 && y_pointer == 48)
||(x_pointer == 36 && y_pointer == 49)
||(x_pointer == 37 && y_pointer == 49)
||(x_pointer == 38 && y_pointer == 49)
||(x_pointer == 39 && y_pointer == 49)
||(x_pointer == 40 && y_pointer == 49)
||(x_pointer == 41 && y_pointer == 49)
||(x_pointer == 42 && y_pointer == 49)
||(x_pointer == 43 && y_pointer == 49)
||(x_pointer == 44 && y_pointer == 49)
||(x_pointer == 45 && y_pointer == 49)
||(x_pointer == 46 && y_pointer == 49)
||(x_pointer == 47 && y_pointer == 49)
||(x_pointer == 48 && y_pointer == 49)
||(x_pointer == 49 && y_pointer == 49)
||(x_pointer == 50 && y_pointer == 49)
||(x_pointer == 51 && y_pointer == 49)
||(x_pointer == 52 && y_pointer == 49)
||(x_pointer == 53 && y_pointer == 49)
||(x_pointer == 54 && y_pointer == 49)
||(x_pointer == 55 && y_pointer == 49)
||(x_pointer == 56 && y_pointer == 49)
||(x_pointer == 57 && y_pointer == 49)
||(x_pointer == 58 && y_pointer == 49)
||(x_pointer == 59 && y_pointer == 49)
||(x_pointer == 60 && y_pointer == 49)
||(x_pointer == 67 && y_pointer == 49)
||(x_pointer == 68 && y_pointer == 49)
||(x_pointer == 69 && y_pointer == 49)
||(x_pointer == 70 && y_pointer == 49)
||(x_pointer == 71 && y_pointer == 49)
||(x_pointer == 72 && y_pointer == 49)
||(x_pointer == 73 && y_pointer == 49)
||(x_pointer == 74 && y_pointer == 49)
||(x_pointer == 75 && y_pointer == 49)
||(x_pointer == 76 && y_pointer == 49)
||(x_pointer == 77 && y_pointer == 49)
||(x_pointer == 78 && y_pointer == 49)
||(x_pointer == 79 && y_pointer == 49)
||(x_pointer == 80 && y_pointer == 49)
||(x_pointer == 81 && y_pointer == 49)
||(x_pointer == 82 && y_pointer == 49)
||(x_pointer == 83 && y_pointer == 49)
||(x_pointer == 84 && y_pointer == 49)
||(x_pointer == 85 && y_pointer == 49)
||(x_pointer == 86 && y_pointer == 49)
||(x_pointer == 87 && y_pointer == 49)
||(x_pointer == 88 && y_pointer == 49)
||(x_pointer == 89 && y_pointer == 49)
||(x_pointer == 96 && y_pointer == 49)
||(x_pointer == 97 && y_pointer == 49)
||(x_pointer == 98 && y_pointer == 49)
||(x_pointer == 99 && y_pointer == 49)
||(x_pointer == 100 && y_pointer == 49)
||(x_pointer == 101 && y_pointer == 49)
||(x_pointer == 102 && y_pointer == 49)
||(x_pointer == 103 && y_pointer == 49)
||(x_pointer == 104 && y_pointer == 49)
||(x_pointer == 105 && y_pointer == 49)
||(x_pointer == 106 && y_pointer == 49)
||(x_pointer == 107 && y_pointer == 49)
||(x_pointer == 108 && y_pointer == 49)
||(x_pointer == 109 && y_pointer == 49)
||(x_pointer == 110 && y_pointer == 49)
||(x_pointer == 111 && y_pointer == 49)
||(x_pointer == 112 && y_pointer == 49)
||(x_pointer == 113 && y_pointer == 49)
||(x_pointer == 114 && y_pointer == 49)
||(x_pointer == 115 && y_pointer == 49)
||(x_pointer == 116 && y_pointer == 49)
||(x_pointer == 117 && y_pointer == 49)
||(x_pointer == 118 && y_pointer == 49)
||(x_pointer == 119 && y_pointer == 49)
||(x_pointer == 120 && y_pointer == 49)
||(x_pointer == 36 && y_pointer == 50)
||(x_pointer == 37 && y_pointer == 50)
||(x_pointer == 38 && y_pointer == 50)
||(x_pointer == 39 && y_pointer == 50)
||(x_pointer == 40 && y_pointer == 50)
||(x_pointer == 41 && y_pointer == 50)
||(x_pointer == 42 && y_pointer == 50)
||(x_pointer == 43 && y_pointer == 50)
||(x_pointer == 44 && y_pointer == 50)
||(x_pointer == 45 && y_pointer == 50)
||(x_pointer == 46 && y_pointer == 50)
||(x_pointer == 47 && y_pointer == 50)
||(x_pointer == 48 && y_pointer == 50)
||(x_pointer == 49 && y_pointer == 50)
||(x_pointer == 50 && y_pointer == 50)
||(x_pointer == 51 && y_pointer == 50)
||(x_pointer == 52 && y_pointer == 50)
||(x_pointer == 53 && y_pointer == 50)
||(x_pointer == 54 && y_pointer == 50)
||(x_pointer == 55 && y_pointer == 50)
||(x_pointer == 56 && y_pointer == 50)
||(x_pointer == 57 && y_pointer == 50)
||(x_pointer == 58 && y_pointer == 50)
||(x_pointer == 59 && y_pointer == 50)
||(x_pointer == 60 && y_pointer == 50)
||(x_pointer == 67 && y_pointer == 50)
||(x_pointer == 68 && y_pointer == 50)
||(x_pointer == 69 && y_pointer == 50)
||(x_pointer == 70 && y_pointer == 50)
||(x_pointer == 71 && y_pointer == 50)
||(x_pointer == 72 && y_pointer == 50)
||(x_pointer == 73 && y_pointer == 50)
||(x_pointer == 74 && y_pointer == 50)
||(x_pointer == 75 && y_pointer == 50)
||(x_pointer == 76 && y_pointer == 50)
||(x_pointer == 77 && y_pointer == 50)
||(x_pointer == 78 && y_pointer == 50)
||(x_pointer == 79 && y_pointer == 50)
||(x_pointer == 80 && y_pointer == 50)
||(x_pointer == 81 && y_pointer == 50)
||(x_pointer == 82 && y_pointer == 50)
||(x_pointer == 83 && y_pointer == 50)
||(x_pointer == 84 && y_pointer == 50)
||(x_pointer == 85 && y_pointer == 50)
||(x_pointer == 86 && y_pointer == 50)
||(x_pointer == 87 && y_pointer == 50)
||(x_pointer == 88 && y_pointer == 50)
||(x_pointer == 89 && y_pointer == 50)
||(x_pointer == 96 && y_pointer == 50)
||(x_pointer == 97 && y_pointer == 50)
||(x_pointer == 98 && y_pointer == 50)
||(x_pointer == 99 && y_pointer == 50)
||(x_pointer == 100 && y_pointer == 50)
||(x_pointer == 101 && y_pointer == 50)
||(x_pointer == 102 && y_pointer == 50)
||(x_pointer == 103 && y_pointer == 50)
||(x_pointer == 104 && y_pointer == 50)
||(x_pointer == 105 && y_pointer == 50)
||(x_pointer == 106 && y_pointer == 50)
||(x_pointer == 107 && y_pointer == 50)
||(x_pointer == 108 && y_pointer == 50)
||(x_pointer == 109 && y_pointer == 50)
||(x_pointer == 110 && y_pointer == 50)
||(x_pointer == 111 && y_pointer == 50)
||(x_pointer == 112 && y_pointer == 50)
||(x_pointer == 113 && y_pointer == 50)
||(x_pointer == 114 && y_pointer == 50)
||(x_pointer == 115 && y_pointer == 50)
||(x_pointer == 116 && y_pointer == 50)
||(x_pointer == 117 && y_pointer == 50)
||(x_pointer == 118 && y_pointer == 50)
||(x_pointer == 119 && y_pointer == 50)
||(x_pointer == 120 && y_pointer == 50)
||(x_pointer == 36 && y_pointer == 51)
||(x_pointer == 37 && y_pointer == 51)
||(x_pointer == 38 && y_pointer == 51)
||(x_pointer == 39 && y_pointer == 51)
||(x_pointer == 40 && y_pointer == 51)
||(x_pointer == 41 && y_pointer == 51)
||(x_pointer == 42 && y_pointer == 51)
||(x_pointer == 43 && y_pointer == 51)
||(x_pointer == 44 && y_pointer == 51)
||(x_pointer == 45 && y_pointer == 51)
||(x_pointer == 46 && y_pointer == 51)
||(x_pointer == 47 && y_pointer == 51)
||(x_pointer == 48 && y_pointer == 51)
||(x_pointer == 49 && y_pointer == 51)
||(x_pointer == 50 && y_pointer == 51)
||(x_pointer == 51 && y_pointer == 51)
||(x_pointer == 52 && y_pointer == 51)
||(x_pointer == 53 && y_pointer == 51)
||(x_pointer == 54 && y_pointer == 51)
||(x_pointer == 55 && y_pointer == 51)
||(x_pointer == 56 && y_pointer == 51)
||(x_pointer == 57 && y_pointer == 51)
||(x_pointer == 58 && y_pointer == 51)
||(x_pointer == 59 && y_pointer == 51)
||(x_pointer == 60 && y_pointer == 51)
||(x_pointer == 67 && y_pointer == 51)
||(x_pointer == 68 && y_pointer == 51)
||(x_pointer == 69 && y_pointer == 51)
||(x_pointer == 70 && y_pointer == 51)
||(x_pointer == 71 && y_pointer == 51)
||(x_pointer == 72 && y_pointer == 51)
||(x_pointer == 73 && y_pointer == 51)
||(x_pointer == 74 && y_pointer == 51)
||(x_pointer == 75 && y_pointer == 51)
||(x_pointer == 76 && y_pointer == 51)
||(x_pointer == 77 && y_pointer == 51)
||(x_pointer == 78 && y_pointer == 51)
||(x_pointer == 79 && y_pointer == 51)
||(x_pointer == 80 && y_pointer == 51)
||(x_pointer == 81 && y_pointer == 51)
||(x_pointer == 82 && y_pointer == 51)
||(x_pointer == 83 && y_pointer == 51)
||(x_pointer == 84 && y_pointer == 51)
||(x_pointer == 85 && y_pointer == 51)
||(x_pointer == 86 && y_pointer == 51)
||(x_pointer == 87 && y_pointer == 51)
||(x_pointer == 88 && y_pointer == 51)
||(x_pointer == 89 && y_pointer == 51)
||(x_pointer == 96 && y_pointer == 51)
||(x_pointer == 97 && y_pointer == 51)
||(x_pointer == 98 && y_pointer == 51)
||(x_pointer == 99 && y_pointer == 51)
||(x_pointer == 100 && y_pointer == 51)
||(x_pointer == 101 && y_pointer == 51)
||(x_pointer == 102 && y_pointer == 51)
||(x_pointer == 103 && y_pointer == 51)
||(x_pointer == 104 && y_pointer == 51)
||(x_pointer == 105 && y_pointer == 51)
||(x_pointer == 106 && y_pointer == 51)
||(x_pointer == 107 && y_pointer == 51)
||(x_pointer == 108 && y_pointer == 51)
||(x_pointer == 109 && y_pointer == 51)
||(x_pointer == 110 && y_pointer == 51)
||(x_pointer == 111 && y_pointer == 51)
||(x_pointer == 112 && y_pointer == 51)
||(x_pointer == 113 && y_pointer == 51)
||(x_pointer == 114 && y_pointer == 51)
||(x_pointer == 115 && y_pointer == 51)
||(x_pointer == 116 && y_pointer == 51)
||(x_pointer == 117 && y_pointer == 51)
||(x_pointer == 118 && y_pointer == 51)
||(x_pointer == 119 && y_pointer == 51)
||(x_pointer == 120 && y_pointer == 51)
||(x_pointer == 36 && y_pointer == 52)
||(x_pointer == 37 && y_pointer == 52)
||(x_pointer == 38 && y_pointer == 52)
||(x_pointer == 39 && y_pointer == 52)
||(x_pointer == 40 && y_pointer == 52)
||(x_pointer == 41 && y_pointer == 52)
||(x_pointer == 42 && y_pointer == 52)
||(x_pointer == 43 && y_pointer == 52)
||(x_pointer == 44 && y_pointer == 52)
||(x_pointer == 45 && y_pointer == 52)
||(x_pointer == 46 && y_pointer == 52)
||(x_pointer == 47 && y_pointer == 52)
||(x_pointer == 48 && y_pointer == 52)
||(x_pointer == 49 && y_pointer == 52)
||(x_pointer == 50 && y_pointer == 52)
||(x_pointer == 51 && y_pointer == 52)
||(x_pointer == 52 && y_pointer == 52)
||(x_pointer == 53 && y_pointer == 52)
||(x_pointer == 54 && y_pointer == 52)
||(x_pointer == 55 && y_pointer == 52)
||(x_pointer == 56 && y_pointer == 52)
||(x_pointer == 57 && y_pointer == 52)
||(x_pointer == 58 && y_pointer == 52)
||(x_pointer == 59 && y_pointer == 52)
||(x_pointer == 60 && y_pointer == 52)
||(x_pointer == 67 && y_pointer == 52)
||(x_pointer == 68 && y_pointer == 52)
||(x_pointer == 69 && y_pointer == 52)
||(x_pointer == 70 && y_pointer == 52)
||(x_pointer == 71 && y_pointer == 52)
||(x_pointer == 72 && y_pointer == 52)
||(x_pointer == 73 && y_pointer == 52)
||(x_pointer == 74 && y_pointer == 52)
||(x_pointer == 75 && y_pointer == 52)
||(x_pointer == 76 && y_pointer == 52)
||(x_pointer == 77 && y_pointer == 52)
||(x_pointer == 78 && y_pointer == 52)
||(x_pointer == 79 && y_pointer == 52)
||(x_pointer == 80 && y_pointer == 52)
||(x_pointer == 81 && y_pointer == 52)
||(x_pointer == 82 && y_pointer == 52)
||(x_pointer == 83 && y_pointer == 52)
||(x_pointer == 84 && y_pointer == 52)
||(x_pointer == 85 && y_pointer == 52)
||(x_pointer == 86 && y_pointer == 52)
||(x_pointer == 87 && y_pointer == 52)
||(x_pointer == 88 && y_pointer == 52)
||(x_pointer == 89 && y_pointer == 52)
||(x_pointer == 96 && y_pointer == 52)
||(x_pointer == 97 && y_pointer == 52)
||(x_pointer == 98 && y_pointer == 52)
||(x_pointer == 99 && y_pointer == 52)
||(x_pointer == 100 && y_pointer == 52)
||(x_pointer == 101 && y_pointer == 52)
||(x_pointer == 102 && y_pointer == 52)
||(x_pointer == 103 && y_pointer == 52)
||(x_pointer == 104 && y_pointer == 52)
||(x_pointer == 105 && y_pointer == 52)
||(x_pointer == 106 && y_pointer == 52)
||(x_pointer == 107 && y_pointer == 52)
||(x_pointer == 108 && y_pointer == 52)
||(x_pointer == 109 && y_pointer == 52)
||(x_pointer == 110 && y_pointer == 52)
||(x_pointer == 111 && y_pointer == 52)
||(x_pointer == 112 && y_pointer == 52)
||(x_pointer == 113 && y_pointer == 52)
||(x_pointer == 114 && y_pointer == 52)
||(x_pointer == 115 && y_pointer == 52)
||(x_pointer == 116 && y_pointer == 52)
||(x_pointer == 117 && y_pointer == 52)
||(x_pointer == 118 && y_pointer == 52)
||(x_pointer == 119 && y_pointer == 52)
||(x_pointer == 120 && y_pointer == 52)
||(x_pointer == 36 && y_pointer == 66)
||(x_pointer == 37 && y_pointer == 66)
||(x_pointer == 38 && y_pointer == 66)
||(x_pointer == 39 && y_pointer == 66)
||(x_pointer == 40 && y_pointer == 66)
||(x_pointer == 41 && y_pointer == 66)
||(x_pointer == 42 && y_pointer == 66)
||(x_pointer == 43 && y_pointer == 66)
||(x_pointer == 44 && y_pointer == 66)
||(x_pointer == 45 && y_pointer == 66)
||(x_pointer == 46 && y_pointer == 66)
||(x_pointer == 47 && y_pointer == 66)
||(x_pointer == 48 && y_pointer == 66)
||(x_pointer == 49 && y_pointer == 66)
||(x_pointer == 50 && y_pointer == 66)
||(x_pointer == 51 && y_pointer == 66)
||(x_pointer == 52 && y_pointer == 66)
||(x_pointer == 53 && y_pointer == 66)
||(x_pointer == 54 && y_pointer == 66)
||(x_pointer == 55 && y_pointer == 66)
||(x_pointer == 56 && y_pointer == 66)
||(x_pointer == 57 && y_pointer == 66)
||(x_pointer == 58 && y_pointer == 66)
||(x_pointer == 59 && y_pointer == 66)
||(x_pointer == 60 && y_pointer == 66)
||(x_pointer == 67 && y_pointer == 66)
||(x_pointer == 68 && y_pointer == 66)
||(x_pointer == 69 && y_pointer == 66)
||(x_pointer == 70 && y_pointer == 66)
||(x_pointer == 71 && y_pointer == 66)
||(x_pointer == 72 && y_pointer == 66)
||(x_pointer == 73 && y_pointer == 66)
||(x_pointer == 74 && y_pointer == 66)
||(x_pointer == 75 && y_pointer == 66)
||(x_pointer == 76 && y_pointer == 66)
||(x_pointer == 77 && y_pointer == 66)
||(x_pointer == 78 && y_pointer == 66)
||(x_pointer == 79 && y_pointer == 66)
||(x_pointer == 80 && y_pointer == 66)
||(x_pointer == 81 && y_pointer == 66)
||(x_pointer == 82 && y_pointer == 66)
||(x_pointer == 83 && y_pointer == 66)
||(x_pointer == 84 && y_pointer == 66)
||(x_pointer == 85 && y_pointer == 66)
||(x_pointer == 86 && y_pointer == 66)
||(x_pointer == 87 && y_pointer == 66)
||(x_pointer == 88 && y_pointer == 66)
||(x_pointer == 89 && y_pointer == 66)
||(x_pointer == 96 && y_pointer == 66)
||(x_pointer == 97 && y_pointer == 66)
||(x_pointer == 98 && y_pointer == 66)
||(x_pointer == 99 && y_pointer == 66)
||(x_pointer == 100 && y_pointer == 66)
||(x_pointer == 101 && y_pointer == 66)
||(x_pointer == 102 && y_pointer == 66)
||(x_pointer == 103 && y_pointer == 66)
||(x_pointer == 104 && y_pointer == 66)
||(x_pointer == 105 && y_pointer == 66)
||(x_pointer == 106 && y_pointer == 66)
||(x_pointer == 107 && y_pointer == 66)
||(x_pointer == 108 && y_pointer == 66)
||(x_pointer == 109 && y_pointer == 66)
||(x_pointer == 110 && y_pointer == 66)
||(x_pointer == 111 && y_pointer == 66)
||(x_pointer == 112 && y_pointer == 66)
||(x_pointer == 113 && y_pointer == 66)
||(x_pointer == 114 && y_pointer == 66)
||(x_pointer == 115 && y_pointer == 66)
||(x_pointer == 116 && y_pointer == 66)
||(x_pointer == 117 && y_pointer == 66)
||(x_pointer == 118 && y_pointer == 66)
||(x_pointer == 119 && y_pointer == 66)
||(x_pointer == 120 && y_pointer == 66)
||(x_pointer == 36 && y_pointer == 67)
||(x_pointer == 37 && y_pointer == 67)
||(x_pointer == 38 && y_pointer == 67)
||(x_pointer == 39 && y_pointer == 67)
||(x_pointer == 40 && y_pointer == 67)
||(x_pointer == 41 && y_pointer == 67)
||(x_pointer == 42 && y_pointer == 67)
||(x_pointer == 43 && y_pointer == 67)
||(x_pointer == 44 && y_pointer == 67)
||(x_pointer == 45 && y_pointer == 67)
||(x_pointer == 46 && y_pointer == 67)
||(x_pointer == 47 && y_pointer == 67)
||(x_pointer == 48 && y_pointer == 67)
||(x_pointer == 49 && y_pointer == 67)
||(x_pointer == 50 && y_pointer == 67)
||(x_pointer == 51 && y_pointer == 67)
||(x_pointer == 52 && y_pointer == 67)
||(x_pointer == 53 && y_pointer == 67)
||(x_pointer == 54 && y_pointer == 67)
||(x_pointer == 55 && y_pointer == 67)
||(x_pointer == 56 && y_pointer == 67)
||(x_pointer == 57 && y_pointer == 67)
||(x_pointer == 58 && y_pointer == 67)
||(x_pointer == 59 && y_pointer == 67)
||(x_pointer == 60 && y_pointer == 67)
||(x_pointer == 67 && y_pointer == 67)
||(x_pointer == 68 && y_pointer == 67)
||(x_pointer == 69 && y_pointer == 67)
||(x_pointer == 70 && y_pointer == 67)
||(x_pointer == 71 && y_pointer == 67)
||(x_pointer == 72 && y_pointer == 67)
||(x_pointer == 73 && y_pointer == 67)
||(x_pointer == 74 && y_pointer == 67)
||(x_pointer == 75 && y_pointer == 67)
||(x_pointer == 76 && y_pointer == 67)
||(x_pointer == 77 && y_pointer == 67)
||(x_pointer == 78 && y_pointer == 67)
||(x_pointer == 79 && y_pointer == 67)
||(x_pointer == 80 && y_pointer == 67)
||(x_pointer == 81 && y_pointer == 67)
||(x_pointer == 82 && y_pointer == 67)
||(x_pointer == 83 && y_pointer == 67)
||(x_pointer == 84 && y_pointer == 67)
||(x_pointer == 85 && y_pointer == 67)
||(x_pointer == 86 && y_pointer == 67)
||(x_pointer == 87 && y_pointer == 67)
||(x_pointer == 88 && y_pointer == 67)
||(x_pointer == 89 && y_pointer == 67)
||(x_pointer == 96 && y_pointer == 67)
||(x_pointer == 97 && y_pointer == 67)
||(x_pointer == 98 && y_pointer == 67)
||(x_pointer == 99 && y_pointer == 67)
||(x_pointer == 100 && y_pointer == 67)
||(x_pointer == 101 && y_pointer == 67)
||(x_pointer == 102 && y_pointer == 67)
||(x_pointer == 103 && y_pointer == 67)
||(x_pointer == 104 && y_pointer == 67)
||(x_pointer == 105 && y_pointer == 67)
||(x_pointer == 106 && y_pointer == 67)
||(x_pointer == 107 && y_pointer == 67)
||(x_pointer == 108 && y_pointer == 67)
||(x_pointer == 109 && y_pointer == 67)
||(x_pointer == 110 && y_pointer == 67)
||(x_pointer == 111 && y_pointer == 67)
||(x_pointer == 112 && y_pointer == 67)
||(x_pointer == 113 && y_pointer == 67)
||(x_pointer == 114 && y_pointer == 67)
||(x_pointer == 115 && y_pointer == 67)
||(x_pointer == 116 && y_pointer == 67)
||(x_pointer == 117 && y_pointer == 67)
||(x_pointer == 118 && y_pointer == 67)
||(x_pointer == 119 && y_pointer == 67)
||(x_pointer == 120 && y_pointer == 67)
||(x_pointer == 36 && y_pointer == 68)
||(x_pointer == 37 && y_pointer == 68)
||(x_pointer == 38 && y_pointer == 68)
||(x_pointer == 39 && y_pointer == 68)
||(x_pointer == 40 && y_pointer == 68)
||(x_pointer == 41 && y_pointer == 68)
||(x_pointer == 42 && y_pointer == 68)
||(x_pointer == 43 && y_pointer == 68)
||(x_pointer == 44 && y_pointer == 68)
||(x_pointer == 45 && y_pointer == 68)
||(x_pointer == 46 && y_pointer == 68)
||(x_pointer == 47 && y_pointer == 68)
||(x_pointer == 48 && y_pointer == 68)
||(x_pointer == 49 && y_pointer == 68)
||(x_pointer == 50 && y_pointer == 68)
||(x_pointer == 51 && y_pointer == 68)
||(x_pointer == 52 && y_pointer == 68)
||(x_pointer == 53 && y_pointer == 68)
||(x_pointer == 54 && y_pointer == 68)
||(x_pointer == 55 && y_pointer == 68)
||(x_pointer == 56 && y_pointer == 68)
||(x_pointer == 57 && y_pointer == 68)
||(x_pointer == 58 && y_pointer == 68)
||(x_pointer == 59 && y_pointer == 68)
||(x_pointer == 60 && y_pointer == 68)
||(x_pointer == 67 && y_pointer == 68)
||(x_pointer == 68 && y_pointer == 68)
||(x_pointer == 69 && y_pointer == 68)
||(x_pointer == 70 && y_pointer == 68)
||(x_pointer == 71 && y_pointer == 68)
||(x_pointer == 72 && y_pointer == 68)
||(x_pointer == 73 && y_pointer == 68)
||(x_pointer == 74 && y_pointer == 68)
||(x_pointer == 75 && y_pointer == 68)
||(x_pointer == 76 && y_pointer == 68)
||(x_pointer == 77 && y_pointer == 68)
||(x_pointer == 78 && y_pointer == 68)
||(x_pointer == 79 && y_pointer == 68)
||(x_pointer == 80 && y_pointer == 68)
||(x_pointer == 81 && y_pointer == 68)
||(x_pointer == 82 && y_pointer == 68)
||(x_pointer == 83 && y_pointer == 68)
||(x_pointer == 84 && y_pointer == 68)
||(x_pointer == 85 && y_pointer == 68)
||(x_pointer == 86 && y_pointer == 68)
||(x_pointer == 87 && y_pointer == 68)
||(x_pointer == 88 && y_pointer == 68)
||(x_pointer == 89 && y_pointer == 68)
||(x_pointer == 96 && y_pointer == 68)
||(x_pointer == 97 && y_pointer == 68)
||(x_pointer == 98 && y_pointer == 68)
||(x_pointer == 99 && y_pointer == 68)
||(x_pointer == 100 && y_pointer == 68)
||(x_pointer == 101 && y_pointer == 68)
||(x_pointer == 102 && y_pointer == 68)
||(x_pointer == 103 && y_pointer == 68)
||(x_pointer == 104 && y_pointer == 68)
||(x_pointer == 105 && y_pointer == 68)
||(x_pointer == 106 && y_pointer == 68)
||(x_pointer == 107 && y_pointer == 68)
||(x_pointer == 108 && y_pointer == 68)
||(x_pointer == 109 && y_pointer == 68)
||(x_pointer == 110 && y_pointer == 68)
||(x_pointer == 111 && y_pointer == 68)
||(x_pointer == 112 && y_pointer == 68)
||(x_pointer == 113 && y_pointer == 68)
||(x_pointer == 114 && y_pointer == 68)
||(x_pointer == 115 && y_pointer == 68)
||(x_pointer == 116 && y_pointer == 68)
||(x_pointer == 117 && y_pointer == 68)
||(x_pointer == 118 && y_pointer == 68)
||(x_pointer == 119 && y_pointer == 68)
||(x_pointer == 120 && y_pointer == 68)
||(x_pointer == 36 && y_pointer == 69)
||(x_pointer == 37 && y_pointer == 69)
||(x_pointer == 38 && y_pointer == 69)
||(x_pointer == 39 && y_pointer == 69)
||(x_pointer == 40 && y_pointer == 69)
||(x_pointer == 41 && y_pointer == 69)
||(x_pointer == 42 && y_pointer == 69)
||(x_pointer == 43 && y_pointer == 69)
||(x_pointer == 44 && y_pointer == 69)
||(x_pointer == 45 && y_pointer == 69)
||(x_pointer == 46 && y_pointer == 69)
||(x_pointer == 47 && y_pointer == 69)
||(x_pointer == 48 && y_pointer == 69)
||(x_pointer == 49 && y_pointer == 69)
||(x_pointer == 50 && y_pointer == 69)
||(x_pointer == 51 && y_pointer == 69)
||(x_pointer == 52 && y_pointer == 69)
||(x_pointer == 53 && y_pointer == 69)
||(x_pointer == 54 && y_pointer == 69)
||(x_pointer == 55 && y_pointer == 69)
||(x_pointer == 56 && y_pointer == 69)
||(x_pointer == 57 && y_pointer == 69)
||(x_pointer == 58 && y_pointer == 69)
||(x_pointer == 59 && y_pointer == 69)
||(x_pointer == 60 && y_pointer == 69)
||(x_pointer == 67 && y_pointer == 69)
||(x_pointer == 68 && y_pointer == 69)
||(x_pointer == 69 && y_pointer == 69)
||(x_pointer == 70 && y_pointer == 69)
||(x_pointer == 71 && y_pointer == 69)
||(x_pointer == 72 && y_pointer == 69)
||(x_pointer == 73 && y_pointer == 69)
||(x_pointer == 74 && y_pointer == 69)
||(x_pointer == 75 && y_pointer == 69)
||(x_pointer == 76 && y_pointer == 69)
||(x_pointer == 77 && y_pointer == 69)
||(x_pointer == 78 && y_pointer == 69)
||(x_pointer == 79 && y_pointer == 69)
||(x_pointer == 80 && y_pointer == 69)
||(x_pointer == 81 && y_pointer == 69)
||(x_pointer == 82 && y_pointer == 69)
||(x_pointer == 83 && y_pointer == 69)
||(x_pointer == 84 && y_pointer == 69)
||(x_pointer == 85 && y_pointer == 69)
||(x_pointer == 86 && y_pointer == 69)
||(x_pointer == 87 && y_pointer == 69)
||(x_pointer == 88 && y_pointer == 69)
||(x_pointer == 89 && y_pointer == 69)
||(x_pointer == 96 && y_pointer == 69)
||(x_pointer == 97 && y_pointer == 69)
||(x_pointer == 98 && y_pointer == 69)
||(x_pointer == 99 && y_pointer == 69)
||(x_pointer == 100 && y_pointer == 69)
||(x_pointer == 101 && y_pointer == 69)
||(x_pointer == 102 && y_pointer == 69)
||(x_pointer == 103 && y_pointer == 69)
||(x_pointer == 104 && y_pointer == 69)
||(x_pointer == 105 && y_pointer == 69)
||(x_pointer == 106 && y_pointer == 69)
||(x_pointer == 107 && y_pointer == 69)
||(x_pointer == 108 && y_pointer == 69)
||(x_pointer == 109 && y_pointer == 69)
||(x_pointer == 110 && y_pointer == 69)
||(x_pointer == 111 && y_pointer == 69)
||(x_pointer == 112 && y_pointer == 69)
||(x_pointer == 113 && y_pointer == 69)
||(x_pointer == 114 && y_pointer == 69)
||(x_pointer == 115 && y_pointer == 69)
||(x_pointer == 116 && y_pointer == 69)
||(x_pointer == 117 && y_pointer == 69)
||(x_pointer == 118 && y_pointer == 69)
||(x_pointer == 119 && y_pointer == 69)
||(x_pointer == 120 && y_pointer == 69)
||(x_pointer == 57 && y_pointer == 70)
||(x_pointer == 58 && y_pointer == 70)
||(x_pointer == 59 && y_pointer == 70)
||(x_pointer == 60 && y_pointer == 70)
||(x_pointer == 67 && y_pointer == 70)
||(x_pointer == 68 && y_pointer == 70)
||(x_pointer == 69 && y_pointer == 70)
||(x_pointer == 70 && y_pointer == 70)
||(x_pointer == 96 && y_pointer == 70)
||(x_pointer == 97 && y_pointer == 70)
||(x_pointer == 98 && y_pointer == 70)
||(x_pointer == 99 && y_pointer == 70)
||(x_pointer == 117 && y_pointer == 70)
||(x_pointer == 118 && y_pointer == 70)
||(x_pointer == 119 && y_pointer == 70)
||(x_pointer == 120 && y_pointer == 70)
||(x_pointer == 57 && y_pointer == 71)
||(x_pointer == 58 && y_pointer == 71)
||(x_pointer == 59 && y_pointer == 71)
||(x_pointer == 60 && y_pointer == 71)
||(x_pointer == 67 && y_pointer == 71)
||(x_pointer == 68 && y_pointer == 71)
||(x_pointer == 69 && y_pointer == 71)
||(x_pointer == 70 && y_pointer == 71)
||(x_pointer == 96 && y_pointer == 71)
||(x_pointer == 97 && y_pointer == 71)
||(x_pointer == 98 && y_pointer == 71)
||(x_pointer == 99 && y_pointer == 71)
||(x_pointer == 117 && y_pointer == 71)
||(x_pointer == 118 && y_pointer == 71)
||(x_pointer == 119 && y_pointer == 71)
||(x_pointer == 120 && y_pointer == 71)
||(x_pointer == 57 && y_pointer == 72)
||(x_pointer == 58 && y_pointer == 72)
||(x_pointer == 59 && y_pointer == 72)
||(x_pointer == 60 && y_pointer == 72)
||(x_pointer == 67 && y_pointer == 72)
||(x_pointer == 68 && y_pointer == 72)
||(x_pointer == 69 && y_pointer == 72)
||(x_pointer == 70 && y_pointer == 72)
||(x_pointer == 96 && y_pointer == 72)
||(x_pointer == 97 && y_pointer == 72)
||(x_pointer == 98 && y_pointer == 72)
||(x_pointer == 99 && y_pointer == 72)
||(x_pointer == 117 && y_pointer == 72)
||(x_pointer == 118 && y_pointer == 72)
||(x_pointer == 119 && y_pointer == 72)
||(x_pointer == 120 && y_pointer == 72)
||(x_pointer == 57 && y_pointer == 73)
||(x_pointer == 58 && y_pointer == 73)
||(x_pointer == 59 && y_pointer == 73)
||(x_pointer == 60 && y_pointer == 73)
||(x_pointer == 67 && y_pointer == 73)
||(x_pointer == 68 && y_pointer == 73)
||(x_pointer == 69 && y_pointer == 73)
||(x_pointer == 70 && y_pointer == 73)
||(x_pointer == 96 && y_pointer == 73)
||(x_pointer == 97 && y_pointer == 73)
||(x_pointer == 98 && y_pointer == 73)
||(x_pointer == 99 && y_pointer == 73)
||(x_pointer == 117 && y_pointer == 73)
||(x_pointer == 118 && y_pointer == 73)
||(x_pointer == 119 && y_pointer == 73)
||(x_pointer == 120 && y_pointer == 73)
||(x_pointer == 57 && y_pointer == 74)
||(x_pointer == 58 && y_pointer == 74)
||(x_pointer == 59 && y_pointer == 74)
||(x_pointer == 60 && y_pointer == 74)
||(x_pointer == 67 && y_pointer == 74)
||(x_pointer == 68 && y_pointer == 74)
||(x_pointer == 69 && y_pointer == 74)
||(x_pointer == 70 && y_pointer == 74)
||(x_pointer == 96 && y_pointer == 74)
||(x_pointer == 97 && y_pointer == 74)
||(x_pointer == 98 && y_pointer == 74)
||(x_pointer == 99 && y_pointer == 74)
||(x_pointer == 117 && y_pointer == 74)
||(x_pointer == 118 && y_pointer == 74)
||(x_pointer == 119 && y_pointer == 74)
||(x_pointer == 120 && y_pointer == 74)
||(x_pointer == 57 && y_pointer == 75)
||(x_pointer == 58 && y_pointer == 75)
||(x_pointer == 59 && y_pointer == 75)
||(x_pointer == 60 && y_pointer == 75)
||(x_pointer == 67 && y_pointer == 75)
||(x_pointer == 68 && y_pointer == 75)
||(x_pointer == 69 && y_pointer == 75)
||(x_pointer == 70 && y_pointer == 75)
||(x_pointer == 96 && y_pointer == 75)
||(x_pointer == 97 && y_pointer == 75)
||(x_pointer == 98 && y_pointer == 75)
||(x_pointer == 99 && y_pointer == 75)
||(x_pointer == 117 && y_pointer == 75)
||(x_pointer == 118 && y_pointer == 75)
||(x_pointer == 119 && y_pointer == 75)
||(x_pointer == 120 && y_pointer == 75)
||(x_pointer == 57 && y_pointer == 76)
||(x_pointer == 58 && y_pointer == 76)
||(x_pointer == 59 && y_pointer == 76)
||(x_pointer == 60 && y_pointer == 76)
||(x_pointer == 67 && y_pointer == 76)
||(x_pointer == 68 && y_pointer == 76)
||(x_pointer == 69 && y_pointer == 76)
||(x_pointer == 70 && y_pointer == 76)
||(x_pointer == 96 && y_pointer == 76)
||(x_pointer == 97 && y_pointer == 76)
||(x_pointer == 98 && y_pointer == 76)
||(x_pointer == 99 && y_pointer == 76)
||(x_pointer == 117 && y_pointer == 76)
||(x_pointer == 118 && y_pointer == 76)
||(x_pointer == 119 && y_pointer == 76)
||(x_pointer == 120 && y_pointer == 76)
||(x_pointer == 57 && y_pointer == 77)
||(x_pointer == 58 && y_pointer == 77)
||(x_pointer == 59 && y_pointer == 77)
||(x_pointer == 60 && y_pointer == 77)
||(x_pointer == 67 && y_pointer == 77)
||(x_pointer == 68 && y_pointer == 77)
||(x_pointer == 69 && y_pointer == 77)
||(x_pointer == 70 && y_pointer == 77)
||(x_pointer == 96 && y_pointer == 77)
||(x_pointer == 97 && y_pointer == 77)
||(x_pointer == 98 && y_pointer == 77)
||(x_pointer == 99 && y_pointer == 77)
||(x_pointer == 117 && y_pointer == 77)
||(x_pointer == 118 && y_pointer == 77)
||(x_pointer == 119 && y_pointer == 77)
||(x_pointer == 120 && y_pointer == 77)
||(x_pointer == 57 && y_pointer == 78)
||(x_pointer == 58 && y_pointer == 78)
||(x_pointer == 59 && y_pointer == 78)
||(x_pointer == 60 && y_pointer == 78)
||(x_pointer == 67 && y_pointer == 78)
||(x_pointer == 68 && y_pointer == 78)
||(x_pointer == 69 && y_pointer == 78)
||(x_pointer == 70 && y_pointer == 78)
||(x_pointer == 96 && y_pointer == 78)
||(x_pointer == 97 && y_pointer == 78)
||(x_pointer == 98 && y_pointer == 78)
||(x_pointer == 99 && y_pointer == 78)
||(x_pointer == 117 && y_pointer == 78)
||(x_pointer == 118 && y_pointer == 78)
||(x_pointer == 119 && y_pointer == 78)
||(x_pointer == 120 && y_pointer == 78)
||(x_pointer == 57 && y_pointer == 79)
||(x_pointer == 58 && y_pointer == 79)
||(x_pointer == 59 && y_pointer == 79)
||(x_pointer == 60 && y_pointer == 79)
||(x_pointer == 67 && y_pointer == 79)
||(x_pointer == 68 && y_pointer == 79)
||(x_pointer == 69 && y_pointer == 79)
||(x_pointer == 70 && y_pointer == 79)
||(x_pointer == 96 && y_pointer == 79)
||(x_pointer == 97 && y_pointer == 79)
||(x_pointer == 98 && y_pointer == 79)
||(x_pointer == 99 && y_pointer == 79)
||(x_pointer == 117 && y_pointer == 79)
||(x_pointer == 118 && y_pointer == 79)
||(x_pointer == 119 && y_pointer == 79)
||(x_pointer == 120 && y_pointer == 79)
||(x_pointer == 36 && y_pointer == 80)
||(x_pointer == 37 && y_pointer == 80)
||(x_pointer == 38 && y_pointer == 80)
||(x_pointer == 39 && y_pointer == 80)
||(x_pointer == 40 && y_pointer == 80)
||(x_pointer == 41 && y_pointer == 80)
||(x_pointer == 42 && y_pointer == 80)
||(x_pointer == 43 && y_pointer == 80)
||(x_pointer == 44 && y_pointer == 80)
||(x_pointer == 45 && y_pointer == 80)
||(x_pointer == 46 && y_pointer == 80)
||(x_pointer == 47 && y_pointer == 80)
||(x_pointer == 48 && y_pointer == 80)
||(x_pointer == 49 && y_pointer == 80)
||(x_pointer == 50 && y_pointer == 80)
||(x_pointer == 51 && y_pointer == 80)
||(x_pointer == 52 && y_pointer == 80)
||(x_pointer == 53 && y_pointer == 80)
||(x_pointer == 54 && y_pointer == 80)
||(x_pointer == 55 && y_pointer == 80)
||(x_pointer == 56 && y_pointer == 80)
||(x_pointer == 57 && y_pointer == 80)
||(x_pointer == 58 && y_pointer == 80)
||(x_pointer == 59 && y_pointer == 80)
||(x_pointer == 60 && y_pointer == 80)
||(x_pointer == 67 && y_pointer == 80)
||(x_pointer == 68 && y_pointer == 80)
||(x_pointer == 69 && y_pointer == 80)
||(x_pointer == 70 && y_pointer == 80)
||(x_pointer == 96 && y_pointer == 80)
||(x_pointer == 97 && y_pointer == 80)
||(x_pointer == 98 && y_pointer == 80)
||(x_pointer == 99 && y_pointer == 80)
||(x_pointer == 100 && y_pointer == 80)
||(x_pointer == 101 && y_pointer == 80)
||(x_pointer == 102 && y_pointer == 80)
||(x_pointer == 103 && y_pointer == 80)
||(x_pointer == 104 && y_pointer == 80)
||(x_pointer == 105 && y_pointer == 80)
||(x_pointer == 106 && y_pointer == 80)
||(x_pointer == 107 && y_pointer == 80)
||(x_pointer == 108 && y_pointer == 80)
||(x_pointer == 109 && y_pointer == 80)
||(x_pointer == 110 && y_pointer == 80)
||(x_pointer == 111 && y_pointer == 80)
||(x_pointer == 112 && y_pointer == 80)
||(x_pointer == 113 && y_pointer == 80)
||(x_pointer == 114 && y_pointer == 80)
||(x_pointer == 115 && y_pointer == 80)
||(x_pointer == 116 && y_pointer == 80)
||(x_pointer == 117 && y_pointer == 80)
||(x_pointer == 118 && y_pointer == 80)
||(x_pointer == 119 && y_pointer == 80)
||(x_pointer == 120 && y_pointer == 80)
||(x_pointer == 36 && y_pointer == 81)
||(x_pointer == 37 && y_pointer == 81)
||(x_pointer == 38 && y_pointer == 81)
||(x_pointer == 39 && y_pointer == 81)
||(x_pointer == 40 && y_pointer == 81)
||(x_pointer == 41 && y_pointer == 81)
||(x_pointer == 42 && y_pointer == 81)
||(x_pointer == 43 && y_pointer == 81)
||(x_pointer == 44 && y_pointer == 81)
||(x_pointer == 45 && y_pointer == 81)
||(x_pointer == 46 && y_pointer == 81)
||(x_pointer == 47 && y_pointer == 81)
||(x_pointer == 48 && y_pointer == 81)
||(x_pointer == 49 && y_pointer == 81)
||(x_pointer == 50 && y_pointer == 81)
||(x_pointer == 51 && y_pointer == 81)
||(x_pointer == 52 && y_pointer == 81)
||(x_pointer == 53 && y_pointer == 81)
||(x_pointer == 54 && y_pointer == 81)
||(x_pointer == 55 && y_pointer == 81)
||(x_pointer == 56 && y_pointer == 81)
||(x_pointer == 57 && y_pointer == 81)
||(x_pointer == 58 && y_pointer == 81)
||(x_pointer == 59 && y_pointer == 81)
||(x_pointer == 60 && y_pointer == 81)
||(x_pointer == 67 && y_pointer == 81)
||(x_pointer == 68 && y_pointer == 81)
||(x_pointer == 69 && y_pointer == 81)
||(x_pointer == 70 && y_pointer == 81)
||(x_pointer == 71 && y_pointer == 81)
||(x_pointer == 72 && y_pointer == 81)
||(x_pointer == 73 && y_pointer == 81)
||(x_pointer == 74 && y_pointer == 81)
||(x_pointer == 75 && y_pointer == 81)
||(x_pointer == 76 && y_pointer == 81)
||(x_pointer == 77 && y_pointer == 81)
||(x_pointer == 78 && y_pointer == 81)
||(x_pointer == 79 && y_pointer == 81)
||(x_pointer == 80 && y_pointer == 81)
||(x_pointer == 81 && y_pointer == 81)
||(x_pointer == 82 && y_pointer == 81)
||(x_pointer == 83 && y_pointer == 81)
||(x_pointer == 84 && y_pointer == 81)
||(x_pointer == 85 && y_pointer == 81)
||(x_pointer == 86 && y_pointer == 81)
||(x_pointer == 87 && y_pointer == 81)
||(x_pointer == 88 && y_pointer == 81)
||(x_pointer == 89 && y_pointer == 81)
||(x_pointer == 96 && y_pointer == 81)
||(x_pointer == 97 && y_pointer == 81)
||(x_pointer == 98 && y_pointer == 81)
||(x_pointer == 99 && y_pointer == 81)
||(x_pointer == 100 && y_pointer == 81)
||(x_pointer == 101 && y_pointer == 81)
||(x_pointer == 102 && y_pointer == 81)
||(x_pointer == 103 && y_pointer == 81)
||(x_pointer == 104 && y_pointer == 81)
||(x_pointer == 105 && y_pointer == 81)
||(x_pointer == 106 && y_pointer == 81)
||(x_pointer == 107 && y_pointer == 81)
||(x_pointer == 108 && y_pointer == 81)
||(x_pointer == 109 && y_pointer == 81)
||(x_pointer == 110 && y_pointer == 81)
||(x_pointer == 111 && y_pointer == 81)
||(x_pointer == 112 && y_pointer == 81)
||(x_pointer == 113 && y_pointer == 81)
||(x_pointer == 114 && y_pointer == 81)
||(x_pointer == 115 && y_pointer == 81)
||(x_pointer == 116 && y_pointer == 81)
||(x_pointer == 117 && y_pointer == 81)
||(x_pointer == 118 && y_pointer == 81)
||(x_pointer == 119 && y_pointer == 81)
||(x_pointer == 120 && y_pointer == 81)
||(x_pointer == 36 && y_pointer == 82)
||(x_pointer == 37 && y_pointer == 82)
||(x_pointer == 38 && y_pointer == 82)
||(x_pointer == 39 && y_pointer == 82)
||(x_pointer == 40 && y_pointer == 82)
||(x_pointer == 41 && y_pointer == 82)
||(x_pointer == 42 && y_pointer == 82)
||(x_pointer == 43 && y_pointer == 82)
||(x_pointer == 44 && y_pointer == 82)
||(x_pointer == 45 && y_pointer == 82)
||(x_pointer == 46 && y_pointer == 82)
||(x_pointer == 47 && y_pointer == 82)
||(x_pointer == 48 && y_pointer == 82)
||(x_pointer == 49 && y_pointer == 82)
||(x_pointer == 50 && y_pointer == 82)
||(x_pointer == 51 && y_pointer == 82)
||(x_pointer == 52 && y_pointer == 82)
||(x_pointer == 53 && y_pointer == 82)
||(x_pointer == 54 && y_pointer == 82)
||(x_pointer == 55 && y_pointer == 82)
||(x_pointer == 56 && y_pointer == 82)
||(x_pointer == 57 && y_pointer == 82)
||(x_pointer == 58 && y_pointer == 82)
||(x_pointer == 59 && y_pointer == 82)
||(x_pointer == 60 && y_pointer == 82)
||(x_pointer == 67 && y_pointer == 82)
||(x_pointer == 68 && y_pointer == 82)
||(x_pointer == 69 && y_pointer == 82)
||(x_pointer == 70 && y_pointer == 82)
||(x_pointer == 71 && y_pointer == 82)
||(x_pointer == 72 && y_pointer == 82)
||(x_pointer == 73 && y_pointer == 82)
||(x_pointer == 74 && y_pointer == 82)
||(x_pointer == 75 && y_pointer == 82)
||(x_pointer == 76 && y_pointer == 82)
||(x_pointer == 77 && y_pointer == 82)
||(x_pointer == 78 && y_pointer == 82)
||(x_pointer == 79 && y_pointer == 82)
||(x_pointer == 80 && y_pointer == 82)
||(x_pointer == 81 && y_pointer == 82)
||(x_pointer == 82 && y_pointer == 82)
||(x_pointer == 83 && y_pointer == 82)
||(x_pointer == 84 && y_pointer == 82)
||(x_pointer == 85 && y_pointer == 82)
||(x_pointer == 86 && y_pointer == 82)
||(x_pointer == 87 && y_pointer == 82)
||(x_pointer == 88 && y_pointer == 82)
||(x_pointer == 89 && y_pointer == 82)
||(x_pointer == 96 && y_pointer == 82)
||(x_pointer == 97 && y_pointer == 82)
||(x_pointer == 98 && y_pointer == 82)
||(x_pointer == 99 && y_pointer == 82)
||(x_pointer == 100 && y_pointer == 82)
||(x_pointer == 101 && y_pointer == 82)
||(x_pointer == 102 && y_pointer == 82)
||(x_pointer == 103 && y_pointer == 82)
||(x_pointer == 104 && y_pointer == 82)
||(x_pointer == 105 && y_pointer == 82)
||(x_pointer == 106 && y_pointer == 82)
||(x_pointer == 107 && y_pointer == 82)
||(x_pointer == 108 && y_pointer == 82)
||(x_pointer == 109 && y_pointer == 82)
||(x_pointer == 110 && y_pointer == 82)
||(x_pointer == 111 && y_pointer == 82)
||(x_pointer == 112 && y_pointer == 82)
||(x_pointer == 113 && y_pointer == 82)
||(x_pointer == 114 && y_pointer == 82)
||(x_pointer == 115 && y_pointer == 82)
||(x_pointer == 116 && y_pointer == 82)
||(x_pointer == 117 && y_pointer == 82)
||(x_pointer == 118 && y_pointer == 82)
||(x_pointer == 119 && y_pointer == 82)
||(x_pointer == 120 && y_pointer == 82)
||(x_pointer == 36 && y_pointer == 83)
||(x_pointer == 37 && y_pointer == 83)
||(x_pointer == 38 && y_pointer == 83)
||(x_pointer == 39 && y_pointer == 83)
||(x_pointer == 40 && y_pointer == 83)
||(x_pointer == 41 && y_pointer == 83)
||(x_pointer == 42 && y_pointer == 83)
||(x_pointer == 43 && y_pointer == 83)
||(x_pointer == 44 && y_pointer == 83)
||(x_pointer == 45 && y_pointer == 83)
||(x_pointer == 46 && y_pointer == 83)
||(x_pointer == 47 && y_pointer == 83)
||(x_pointer == 48 && y_pointer == 83)
||(x_pointer == 49 && y_pointer == 83)
||(x_pointer == 50 && y_pointer == 83)
||(x_pointer == 51 && y_pointer == 83)
||(x_pointer == 52 && y_pointer == 83)
||(x_pointer == 53 && y_pointer == 83)
||(x_pointer == 54 && y_pointer == 83)
||(x_pointer == 55 && y_pointer == 83)
||(x_pointer == 56 && y_pointer == 83)
||(x_pointer == 57 && y_pointer == 83)
||(x_pointer == 58 && y_pointer == 83)
||(x_pointer == 59 && y_pointer == 83)
||(x_pointer == 60 && y_pointer == 83)
||(x_pointer == 67 && y_pointer == 83)
||(x_pointer == 68 && y_pointer == 83)
||(x_pointer == 69 && y_pointer == 83)
||(x_pointer == 70 && y_pointer == 83)
||(x_pointer == 71 && y_pointer == 83)
||(x_pointer == 72 && y_pointer == 83)
||(x_pointer == 73 && y_pointer == 83)
||(x_pointer == 74 && y_pointer == 83)
||(x_pointer == 75 && y_pointer == 83)
||(x_pointer == 76 && y_pointer == 83)
||(x_pointer == 77 && y_pointer == 83)
||(x_pointer == 78 && y_pointer == 83)
||(x_pointer == 79 && y_pointer == 83)
||(x_pointer == 80 && y_pointer == 83)
||(x_pointer == 81 && y_pointer == 83)
||(x_pointer == 82 && y_pointer == 83)
||(x_pointer == 83 && y_pointer == 83)
||(x_pointer == 84 && y_pointer == 83)
||(x_pointer == 85 && y_pointer == 83)
||(x_pointer == 86 && y_pointer == 83)
||(x_pointer == 87 && y_pointer == 83)
||(x_pointer == 88 && y_pointer == 83)
||(x_pointer == 89 && y_pointer == 83)
||(x_pointer == 96 && y_pointer == 83)
||(x_pointer == 97 && y_pointer == 83)
||(x_pointer == 98 && y_pointer == 83)
||(x_pointer == 99 && y_pointer == 83)
||(x_pointer == 100 && y_pointer == 83)
||(x_pointer == 101 && y_pointer == 83)
||(x_pointer == 102 && y_pointer == 83)
||(x_pointer == 103 && y_pointer == 83)
||(x_pointer == 104 && y_pointer == 83)
||(x_pointer == 105 && y_pointer == 83)
||(x_pointer == 106 && y_pointer == 83)
||(x_pointer == 107 && y_pointer == 83)
||(x_pointer == 108 && y_pointer == 83)
||(x_pointer == 109 && y_pointer == 83)
||(x_pointer == 110 && y_pointer == 83)
||(x_pointer == 111 && y_pointer == 83)
||(x_pointer == 112 && y_pointer == 83)
||(x_pointer == 113 && y_pointer == 83)
||(x_pointer == 114 && y_pointer == 83)
||(x_pointer == 115 && y_pointer == 83)
||(x_pointer == 116 && y_pointer == 83)
||(x_pointer == 117 && y_pointer == 83)
||(x_pointer == 118 && y_pointer == 83)
||(x_pointer == 119 && y_pointer == 83)
||(x_pointer == 120 && y_pointer == 83)
||(x_pointer == 36 && y_pointer == 84)
||(x_pointer == 37 && y_pointer == 84)
||(x_pointer == 38 && y_pointer == 84)
||(x_pointer == 39 && y_pointer == 84)
||(x_pointer == 67 && y_pointer == 84)
||(x_pointer == 68 && y_pointer == 84)
||(x_pointer == 69 && y_pointer == 84)
||(x_pointer == 70 && y_pointer == 84)
||(x_pointer == 71 && y_pointer == 84)
||(x_pointer == 72 && y_pointer == 84)
||(x_pointer == 73 && y_pointer == 84)
||(x_pointer == 74 && y_pointer == 84)
||(x_pointer == 75 && y_pointer == 84)
||(x_pointer == 76 && y_pointer == 84)
||(x_pointer == 77 && y_pointer == 84)
||(x_pointer == 78 && y_pointer == 84)
||(x_pointer == 79 && y_pointer == 84)
||(x_pointer == 80 && y_pointer == 84)
||(x_pointer == 81 && y_pointer == 84)
||(x_pointer == 82 && y_pointer == 84)
||(x_pointer == 83 && y_pointer == 84)
||(x_pointer == 84 && y_pointer == 84)
||(x_pointer == 85 && y_pointer == 84)
||(x_pointer == 86 && y_pointer == 84)
||(x_pointer == 87 && y_pointer == 84)
||(x_pointer == 88 && y_pointer == 84)
||(x_pointer == 89 && y_pointer == 84)
||(x_pointer == 96 && y_pointer == 84)
||(x_pointer == 97 && y_pointer == 84)
||(x_pointer == 98 && y_pointer == 84)
||(x_pointer == 99 && y_pointer == 84)
||(x_pointer == 100 && y_pointer == 84)
||(x_pointer == 101 && y_pointer == 84)
||(x_pointer == 102 && y_pointer == 84)
||(x_pointer == 103 && y_pointer == 84)
||(x_pointer == 104 && y_pointer == 84)
||(x_pointer == 105 && y_pointer == 84)
||(x_pointer == 106 && y_pointer == 84)
||(x_pointer == 107 && y_pointer == 84)
||(x_pointer == 108 && y_pointer == 84)
||(x_pointer == 109 && y_pointer == 84)
||(x_pointer == 110 && y_pointer == 84)
||(x_pointer == 111 && y_pointer == 84)
||(x_pointer == 112 && y_pointer == 84)
||(x_pointer == 113 && y_pointer == 84)
||(x_pointer == 114 && y_pointer == 84)
||(x_pointer == 115 && y_pointer == 84)
||(x_pointer == 116 && y_pointer == 84)
||(x_pointer == 117 && y_pointer == 84)
||(x_pointer == 118 && y_pointer == 84)
||(x_pointer == 119 && y_pointer == 84)
||(x_pointer == 120 && y_pointer == 84)
||(x_pointer == 36 && y_pointer == 85)
||(x_pointer == 37 && y_pointer == 85)
||(x_pointer == 38 && y_pointer == 85)
||(x_pointer == 39 && y_pointer == 85)
||(x_pointer == 86 && y_pointer == 85)
||(x_pointer == 87 && y_pointer == 85)
||(x_pointer == 88 && y_pointer == 85)
||(x_pointer == 89 && y_pointer == 85)
||(x_pointer == 96 && y_pointer == 85)
||(x_pointer == 97 && y_pointer == 85)
||(x_pointer == 98 && y_pointer == 85)
||(x_pointer == 99 && y_pointer == 85)
||(x_pointer == 117 && y_pointer == 85)
||(x_pointer == 118 && y_pointer == 85)
||(x_pointer == 119 && y_pointer == 85)
||(x_pointer == 120 && y_pointer == 85)
||(x_pointer == 36 && y_pointer == 86)
||(x_pointer == 37 && y_pointer == 86)
||(x_pointer == 38 && y_pointer == 86)
||(x_pointer == 39 && y_pointer == 86)
||(x_pointer == 86 && y_pointer == 86)
||(x_pointer == 87 && y_pointer == 86)
||(x_pointer == 88 && y_pointer == 86)
||(x_pointer == 89 && y_pointer == 86)
||(x_pointer == 96 && y_pointer == 86)
||(x_pointer == 97 && y_pointer == 86)
||(x_pointer == 98 && y_pointer == 86)
||(x_pointer == 99 && y_pointer == 86)
||(x_pointer == 117 && y_pointer == 86)
||(x_pointer == 118 && y_pointer == 86)
||(x_pointer == 119 && y_pointer == 86)
||(x_pointer == 120 && y_pointer == 86)
||(x_pointer == 36 && y_pointer == 87)
||(x_pointer == 37 && y_pointer == 87)
||(x_pointer == 38 && y_pointer == 87)
||(x_pointer == 39 && y_pointer == 87)
||(x_pointer == 86 && y_pointer == 87)
||(x_pointer == 87 && y_pointer == 87)
||(x_pointer == 88 && y_pointer == 87)
||(x_pointer == 89 && y_pointer == 87)
||(x_pointer == 96 && y_pointer == 87)
||(x_pointer == 97 && y_pointer == 87)
||(x_pointer == 98 && y_pointer == 87)
||(x_pointer == 99 && y_pointer == 87)
||(x_pointer == 117 && y_pointer == 87)
||(x_pointer == 118 && y_pointer == 87)
||(x_pointer == 119 && y_pointer == 87)
||(x_pointer == 120 && y_pointer == 87)
||(x_pointer == 36 && y_pointer == 88)
||(x_pointer == 37 && y_pointer == 88)
||(x_pointer == 38 && y_pointer == 88)
||(x_pointer == 39 && y_pointer == 88)
||(x_pointer == 86 && y_pointer == 88)
||(x_pointer == 87 && y_pointer == 88)
||(x_pointer == 88 && y_pointer == 88)
||(x_pointer == 89 && y_pointer == 88)
||(x_pointer == 96 && y_pointer == 88)
||(x_pointer == 97 && y_pointer == 88)
||(x_pointer == 98 && y_pointer == 88)
||(x_pointer == 99 && y_pointer == 88)
||(x_pointer == 117 && y_pointer == 88)
||(x_pointer == 118 && y_pointer == 88)
||(x_pointer == 119 && y_pointer == 88)
||(x_pointer == 120 && y_pointer == 88)
||(x_pointer == 36 && y_pointer == 89)
||(x_pointer == 37 && y_pointer == 89)
||(x_pointer == 38 && y_pointer == 89)
||(x_pointer == 39 && y_pointer == 89)
||(x_pointer == 86 && y_pointer == 89)
||(x_pointer == 87 && y_pointer == 89)
||(x_pointer == 88 && y_pointer == 89)
||(x_pointer == 89 && y_pointer == 89)
||(x_pointer == 96 && y_pointer == 89)
||(x_pointer == 97 && y_pointer == 89)
||(x_pointer == 98 && y_pointer == 89)
||(x_pointer == 99 && y_pointer == 89)
||(x_pointer == 117 && y_pointer == 89)
||(x_pointer == 118 && y_pointer == 89)
||(x_pointer == 119 && y_pointer == 89)
||(x_pointer == 120 && y_pointer == 89)
||(x_pointer == 36 && y_pointer == 90)
||(x_pointer == 37 && y_pointer == 90)
||(x_pointer == 38 && y_pointer == 90)
||(x_pointer == 39 && y_pointer == 90)
||(x_pointer == 86 && y_pointer == 90)
||(x_pointer == 87 && y_pointer == 90)
||(x_pointer == 88 && y_pointer == 90)
||(x_pointer == 89 && y_pointer == 90)
||(x_pointer == 96 && y_pointer == 90)
||(x_pointer == 97 && y_pointer == 90)
||(x_pointer == 98 && y_pointer == 90)
||(x_pointer == 99 && y_pointer == 90)
||(x_pointer == 117 && y_pointer == 90)
||(x_pointer == 118 && y_pointer == 90)
||(x_pointer == 119 && y_pointer == 90)
||(x_pointer == 120 && y_pointer == 90)
||(x_pointer == 36 && y_pointer == 91)
||(x_pointer == 37 && y_pointer == 91)
||(x_pointer == 38 && y_pointer == 91)
||(x_pointer == 39 && y_pointer == 91)
||(x_pointer == 86 && y_pointer == 91)
||(x_pointer == 87 && y_pointer == 91)
||(x_pointer == 88 && y_pointer == 91)
||(x_pointer == 89 && y_pointer == 91)
||(x_pointer == 96 && y_pointer == 91)
||(x_pointer == 97 && y_pointer == 91)
||(x_pointer == 98 && y_pointer == 91)
||(x_pointer == 99 && y_pointer == 91)
||(x_pointer == 117 && y_pointer == 91)
||(x_pointer == 118 && y_pointer == 91)
||(x_pointer == 119 && y_pointer == 91)
||(x_pointer == 120 && y_pointer == 91)
||(x_pointer == 36 && y_pointer == 92)
||(x_pointer == 37 && y_pointer == 92)
||(x_pointer == 38 && y_pointer == 92)
||(x_pointer == 39 && y_pointer == 92)
||(x_pointer == 86 && y_pointer == 92)
||(x_pointer == 87 && y_pointer == 92)
||(x_pointer == 88 && y_pointer == 92)
||(x_pointer == 89 && y_pointer == 92)
||(x_pointer == 96 && y_pointer == 92)
||(x_pointer == 97 && y_pointer == 92)
||(x_pointer == 98 && y_pointer == 92)
||(x_pointer == 99 && y_pointer == 92)
||(x_pointer == 117 && y_pointer == 92)
||(x_pointer == 118 && y_pointer == 92)
||(x_pointer == 119 && y_pointer == 92)
||(x_pointer == 120 && y_pointer == 92)
||(x_pointer == 36 && y_pointer == 93)
||(x_pointer == 37 && y_pointer == 93)
||(x_pointer == 38 && y_pointer == 93)
||(x_pointer == 39 && y_pointer == 93)
||(x_pointer == 86 && y_pointer == 93)
||(x_pointer == 87 && y_pointer == 93)
||(x_pointer == 88 && y_pointer == 93)
||(x_pointer == 89 && y_pointer == 93)
||(x_pointer == 96 && y_pointer == 93)
||(x_pointer == 97 && y_pointer == 93)
||(x_pointer == 98 && y_pointer == 93)
||(x_pointer == 99 && y_pointer == 93)
||(x_pointer == 117 && y_pointer == 93)
||(x_pointer == 118 && y_pointer == 93)
||(x_pointer == 119 && y_pointer == 93)
||(x_pointer == 120 && y_pointer == 93)
||(x_pointer == 36 && y_pointer == 94)
||(x_pointer == 37 && y_pointer == 94)
||(x_pointer == 38 && y_pointer == 94)
||(x_pointer == 39 && y_pointer == 94)
||(x_pointer == 40 && y_pointer == 94)
||(x_pointer == 41 && y_pointer == 94)
||(x_pointer == 42 && y_pointer == 94)
||(x_pointer == 43 && y_pointer == 94)
||(x_pointer == 44 && y_pointer == 94)
||(x_pointer == 45 && y_pointer == 94)
||(x_pointer == 46 && y_pointer == 94)
||(x_pointer == 47 && y_pointer == 94)
||(x_pointer == 48 && y_pointer == 94)
||(x_pointer == 49 && y_pointer == 94)
||(x_pointer == 50 && y_pointer == 94)
||(x_pointer == 51 && y_pointer == 94)
||(x_pointer == 52 && y_pointer == 94)
||(x_pointer == 53 && y_pointer == 94)
||(x_pointer == 54 && y_pointer == 94)
||(x_pointer == 55 && y_pointer == 94)
||(x_pointer == 56 && y_pointer == 94)
||(x_pointer == 57 && y_pointer == 94)
||(x_pointer == 58 && y_pointer == 94)
||(x_pointer == 59 && y_pointer == 94)
||(x_pointer == 60 && y_pointer == 94)
||(x_pointer == 67 && y_pointer == 94)
||(x_pointer == 68 && y_pointer == 94)
||(x_pointer == 69 && y_pointer == 94)
||(x_pointer == 70 && y_pointer == 94)
||(x_pointer == 71 && y_pointer == 94)
||(x_pointer == 72 && y_pointer == 94)
||(x_pointer == 73 && y_pointer == 94)
||(x_pointer == 74 && y_pointer == 94)
||(x_pointer == 75 && y_pointer == 94)
||(x_pointer == 76 && y_pointer == 94)
||(x_pointer == 77 && y_pointer == 94)
||(x_pointer == 78 && y_pointer == 94)
||(x_pointer == 79 && y_pointer == 94)
||(x_pointer == 80 && y_pointer == 94)
||(x_pointer == 81 && y_pointer == 94)
||(x_pointer == 82 && y_pointer == 94)
||(x_pointer == 83 && y_pointer == 94)
||(x_pointer == 84 && y_pointer == 94)
||(x_pointer == 85 && y_pointer == 94)
||(x_pointer == 86 && y_pointer == 94)
||(x_pointer == 87 && y_pointer == 94)
||(x_pointer == 88 && y_pointer == 94)
||(x_pointer == 89 && y_pointer == 94)
||(x_pointer == 96 && y_pointer == 94)
||(x_pointer == 97 && y_pointer == 94)
||(x_pointer == 98 && y_pointer == 94)
||(x_pointer == 99 && y_pointer == 94)
||(x_pointer == 100 && y_pointer == 94)
||(x_pointer == 101 && y_pointer == 94)
||(x_pointer == 102 && y_pointer == 94)
||(x_pointer == 103 && y_pointer == 94)
||(x_pointer == 104 && y_pointer == 94)
||(x_pointer == 105 && y_pointer == 94)
||(x_pointer == 106 && y_pointer == 94)
||(x_pointer == 107 && y_pointer == 94)
||(x_pointer == 108 && y_pointer == 94)
||(x_pointer == 109 && y_pointer == 94)
||(x_pointer == 110 && y_pointer == 94)
||(x_pointer == 111 && y_pointer == 94)
||(x_pointer == 112 && y_pointer == 94)
||(x_pointer == 113 && y_pointer == 94)
||(x_pointer == 114 && y_pointer == 94)
||(x_pointer == 115 && y_pointer == 94)
||(x_pointer == 116 && y_pointer == 94)
||(x_pointer == 117 && y_pointer == 94)
||(x_pointer == 118 && y_pointer == 94)
||(x_pointer == 119 && y_pointer == 94)
||(x_pointer == 120 && y_pointer == 94)
||(x_pointer == 36 && y_pointer == 95)
||(x_pointer == 37 && y_pointer == 95)
||(x_pointer == 38 && y_pointer == 95)
||(x_pointer == 39 && y_pointer == 95)
||(x_pointer == 40 && y_pointer == 95)
||(x_pointer == 41 && y_pointer == 95)
||(x_pointer == 42 && y_pointer == 95)
||(x_pointer == 43 && y_pointer == 95)
||(x_pointer == 44 && y_pointer == 95)
||(x_pointer == 45 && y_pointer == 95)
||(x_pointer == 46 && y_pointer == 95)
||(x_pointer == 47 && y_pointer == 95)
||(x_pointer == 48 && y_pointer == 95)
||(x_pointer == 49 && y_pointer == 95)
||(x_pointer == 50 && y_pointer == 95)
||(x_pointer == 51 && y_pointer == 95)
||(x_pointer == 52 && y_pointer == 95)
||(x_pointer == 53 && y_pointer == 95)
||(x_pointer == 54 && y_pointer == 95)
||(x_pointer == 55 && y_pointer == 95)
||(x_pointer == 56 && y_pointer == 95)
||(x_pointer == 57 && y_pointer == 95)
||(x_pointer == 58 && y_pointer == 95)
||(x_pointer == 59 && y_pointer == 95)
||(x_pointer == 60 && y_pointer == 95)
||(x_pointer == 67 && y_pointer == 95)
||(x_pointer == 68 && y_pointer == 95)
||(x_pointer == 69 && y_pointer == 95)
||(x_pointer == 70 && y_pointer == 95)
||(x_pointer == 71 && y_pointer == 95)
||(x_pointer == 72 && y_pointer == 95)
||(x_pointer == 73 && y_pointer == 95)
||(x_pointer == 74 && y_pointer == 95)
||(x_pointer == 75 && y_pointer == 95)
||(x_pointer == 76 && y_pointer == 95)
||(x_pointer == 77 && y_pointer == 95)
||(x_pointer == 78 && y_pointer == 95)
||(x_pointer == 79 && y_pointer == 95)
||(x_pointer == 80 && y_pointer == 95)
||(x_pointer == 81 && y_pointer == 95)
||(x_pointer == 82 && y_pointer == 95)
||(x_pointer == 83 && y_pointer == 95)
||(x_pointer == 84 && y_pointer == 95)
||(x_pointer == 85 && y_pointer == 95)
||(x_pointer == 86 && y_pointer == 95)
||(x_pointer == 87 && y_pointer == 95)
||(x_pointer == 88 && y_pointer == 95)
||(x_pointer == 89 && y_pointer == 95)
||(x_pointer == 96 && y_pointer == 95)
||(x_pointer == 97 && y_pointer == 95)
||(x_pointer == 98 && y_pointer == 95)
||(x_pointer == 99 && y_pointer == 95)
||(x_pointer == 100 && y_pointer == 95)
||(x_pointer == 101 && y_pointer == 95)
||(x_pointer == 102 && y_pointer == 95)
||(x_pointer == 103 && y_pointer == 95)
||(x_pointer == 104 && y_pointer == 95)
||(x_pointer == 105 && y_pointer == 95)
||(x_pointer == 106 && y_pointer == 95)
||(x_pointer == 107 && y_pointer == 95)
||(x_pointer == 108 && y_pointer == 95)
||(x_pointer == 109 && y_pointer == 95)
||(x_pointer == 110 && y_pointer == 95)
||(x_pointer == 111 && y_pointer == 95)
||(x_pointer == 112 && y_pointer == 95)
||(x_pointer == 113 && y_pointer == 95)
||(x_pointer == 114 && y_pointer == 95)
||(x_pointer == 115 && y_pointer == 95)
||(x_pointer == 116 && y_pointer == 95)
||(x_pointer == 117 && y_pointer == 95)
||(x_pointer == 118 && y_pointer == 95)
||(x_pointer == 119 && y_pointer == 95)
||(x_pointer == 120 && y_pointer == 95)
||(x_pointer == 36 && y_pointer == 96)
||(x_pointer == 37 && y_pointer == 96)
||(x_pointer == 38 && y_pointer == 96)
||(x_pointer == 39 && y_pointer == 96)
||(x_pointer == 40 && y_pointer == 96)
||(x_pointer == 41 && y_pointer == 96)
||(x_pointer == 42 && y_pointer == 96)
||(x_pointer == 43 && y_pointer == 96)
||(x_pointer == 44 && y_pointer == 96)
||(x_pointer == 45 && y_pointer == 96)
||(x_pointer == 46 && y_pointer == 96)
||(x_pointer == 47 && y_pointer == 96)
||(x_pointer == 48 && y_pointer == 96)
||(x_pointer == 49 && y_pointer == 96)
||(x_pointer == 50 && y_pointer == 96)
||(x_pointer == 51 && y_pointer == 96)
||(x_pointer == 52 && y_pointer == 96)
||(x_pointer == 53 && y_pointer == 96)
||(x_pointer == 54 && y_pointer == 96)
||(x_pointer == 55 && y_pointer == 96)
||(x_pointer == 56 && y_pointer == 96)
||(x_pointer == 57 && y_pointer == 96)
||(x_pointer == 58 && y_pointer == 96)
||(x_pointer == 59 && y_pointer == 96)
||(x_pointer == 60 && y_pointer == 96)
||(x_pointer == 67 && y_pointer == 96)
||(x_pointer == 68 && y_pointer == 96)
||(x_pointer == 69 && y_pointer == 96)
||(x_pointer == 70 && y_pointer == 96)
||(x_pointer == 71 && y_pointer == 96)
||(x_pointer == 72 && y_pointer == 96)
||(x_pointer == 73 && y_pointer == 96)
||(x_pointer == 74 && y_pointer == 96)
||(x_pointer == 75 && y_pointer == 96)
||(x_pointer == 76 && y_pointer == 96)
||(x_pointer == 77 && y_pointer == 96)
||(x_pointer == 78 && y_pointer == 96)
||(x_pointer == 79 && y_pointer == 96)
||(x_pointer == 80 && y_pointer == 96)
||(x_pointer == 81 && y_pointer == 96)
||(x_pointer == 82 && y_pointer == 96)
||(x_pointer == 83 && y_pointer == 96)
||(x_pointer == 84 && y_pointer == 96)
||(x_pointer == 85 && y_pointer == 96)
||(x_pointer == 86 && y_pointer == 96)
||(x_pointer == 87 && y_pointer == 96)
||(x_pointer == 88 && y_pointer == 96)
||(x_pointer == 89 && y_pointer == 96)
||(x_pointer == 96 && y_pointer == 96)
||(x_pointer == 97 && y_pointer == 96)
||(x_pointer == 98 && y_pointer == 96)
||(x_pointer == 99 && y_pointer == 96)
||(x_pointer == 100 && y_pointer == 96)
||(x_pointer == 101 && y_pointer == 96)
||(x_pointer == 102 && y_pointer == 96)
||(x_pointer == 103 && y_pointer == 96)
||(x_pointer == 104 && y_pointer == 96)
||(x_pointer == 105 && y_pointer == 96)
||(x_pointer == 106 && y_pointer == 96)
||(x_pointer == 107 && y_pointer == 96)
||(x_pointer == 108 && y_pointer == 96)
||(x_pointer == 109 && y_pointer == 96)
||(x_pointer == 110 && y_pointer == 96)
||(x_pointer == 111 && y_pointer == 96)
||(x_pointer == 112 && y_pointer == 96)
||(x_pointer == 113 && y_pointer == 96)
||(x_pointer == 114 && y_pointer == 96)
||(x_pointer == 115 && y_pointer == 96)
||(x_pointer == 116 && y_pointer == 96)
||(x_pointer == 117 && y_pointer == 96)
||(x_pointer == 118 && y_pointer == 96)
||(x_pointer == 119 && y_pointer == 96)
||(x_pointer == 120 && y_pointer == 96)
||(x_pointer == 36 && y_pointer == 97)
||(x_pointer == 37 && y_pointer == 97)
||(x_pointer == 38 && y_pointer == 97)
||(x_pointer == 39 && y_pointer == 97)
||(x_pointer == 40 && y_pointer == 97)
||(x_pointer == 41 && y_pointer == 97)
||(x_pointer == 42 && y_pointer == 97)
||(x_pointer == 43 && y_pointer == 97)
||(x_pointer == 44 && y_pointer == 97)
||(x_pointer == 45 && y_pointer == 97)
||(x_pointer == 46 && y_pointer == 97)
||(x_pointer == 47 && y_pointer == 97)
||(x_pointer == 48 && y_pointer == 97)
||(x_pointer == 49 && y_pointer == 97)
||(x_pointer == 50 && y_pointer == 97)
||(x_pointer == 51 && y_pointer == 97)
||(x_pointer == 52 && y_pointer == 97)
||(x_pointer == 53 && y_pointer == 97)
||(x_pointer == 54 && y_pointer == 97)
||(x_pointer == 55 && y_pointer == 97)
||(x_pointer == 56 && y_pointer == 97)
||(x_pointer == 57 && y_pointer == 97)
||(x_pointer == 58 && y_pointer == 97)
||(x_pointer == 59 && y_pointer == 97)
||(x_pointer == 60 && y_pointer == 97)
||(x_pointer == 67 && y_pointer == 97)
||(x_pointer == 68 && y_pointer == 97)
||(x_pointer == 69 && y_pointer == 97)
||(x_pointer == 70 && y_pointer == 97)
||(x_pointer == 71 && y_pointer == 97)
||(x_pointer == 72 && y_pointer == 97)
||(x_pointer == 73 && y_pointer == 97)
||(x_pointer == 74 && y_pointer == 97)
||(x_pointer == 75 && y_pointer == 97)
||(x_pointer == 76 && y_pointer == 97)
||(x_pointer == 77 && y_pointer == 97)
||(x_pointer == 78 && y_pointer == 97)
||(x_pointer == 79 && y_pointer == 97)
||(x_pointer == 80 && y_pointer == 97)
||(x_pointer == 81 && y_pointer == 97)
||(x_pointer == 82 && y_pointer == 97)
||(x_pointer == 83 && y_pointer == 97)
||(x_pointer == 84 && y_pointer == 97)
||(x_pointer == 85 && y_pointer == 97)
||(x_pointer == 86 && y_pointer == 97)
||(x_pointer == 87 && y_pointer == 97)
||(x_pointer == 88 && y_pointer == 97)
||(x_pointer == 89 && y_pointer == 97)
||(x_pointer == 96 && y_pointer == 97)
||(x_pointer == 97 && y_pointer == 97)
||(x_pointer == 98 && y_pointer == 97)
||(x_pointer == 99 && y_pointer == 97)
||(x_pointer == 100 && y_pointer == 97)
||(x_pointer == 101 && y_pointer == 97)
||(x_pointer == 102 && y_pointer == 97)
||(x_pointer == 103 && y_pointer == 97)
||(x_pointer == 104 && y_pointer == 97)
||(x_pointer == 105 && y_pointer == 97)
||(x_pointer == 106 && y_pointer == 97)
||(x_pointer == 107 && y_pointer == 97)
||(x_pointer == 108 && y_pointer == 97)
||(x_pointer == 109 && y_pointer == 97)
||(x_pointer == 110 && y_pointer == 97)
||(x_pointer == 111 && y_pointer == 97)
||(x_pointer == 112 && y_pointer == 97)
||(x_pointer == 113 && y_pointer == 97)
||(x_pointer == 114 && y_pointer == 97)
||(x_pointer == 115 && y_pointer == 97)
||(x_pointer == 116 && y_pointer == 97)
||(x_pointer == 117 && y_pointer == 97)
||(x_pointer == 118 && y_pointer == 97)
||(x_pointer == 119 && y_pointer == 97)
||(x_pointer == 120 && y_pointer == 97));
endmodule